PK   ��X7���;!  )?    cirkitFile.json�ݒ�ȑ�_���G4��B$z��Yox"v~bg�� GSd����лo%HI�A��}a�h$��Ï��D��a��~n6�b�kʟ���j���Iv;yS��w��G���~�)���]u�fr�A�����7�|�T�|ǔ�i��l����<	K?K
�IXTռIӺjJW����׷�^AZ�/�۷��M�ٗ��BB!����%!w.���e���|����$�abyqW�_,��ߛ�
�L�V���`Up�2X\���
����
����
�,�V�X����,) U�*)��R��T�����w�Z�A���^��^����^����^����^����^����^��qNg��f�Ha��f�H���뮷Oq���^;���^;���^;���^;���^;�N�Gf
{�L��,)��,)��,) ��3��N�D���N�D���N�D���N�D���N�D���N��+��v�%"��v�%"��v�%"��v�%"�⪽v{�4KD
{�4KD
{�4KD
{�4KD
{�4K�2��N�D���N�D���N�D���N�D���N�D� |5e����v�%"��v�%"��v�%"��v�%\��k�Y"R�k�Y"R�kgG�~���%�j�|OGy�]W���}����4?�K'X:��l�t��s����cc�,�+Sl�Rl�t�������N�tq��]���N�t�l��]���N�t��bc7��J'X:Wΰ��ac�,�+l�
l�t��ӻ��c����	�O���.���/l0�0�|���O���,�����Wp��N�'`>�o?����	�O�8��8�|��{����,����.op����'`>�??����	�O�_`�,���tM 8~`���0��f ���+���`�����'`>]A��`�̧k_���,���t�8~`���0��7��?�|�ӕR�����O�|��?����	�OW��o� �,���t]8~`���0����?�|�ӵ�����B�f�)��`���0����?�|�ӕ������O�|�f?����	�OW���X>��:ip����'`>]ፍ_ �,���tm:8~`���0�����?�|��~ �����O�|�� ?�J�R��`����'`>���`�̧}/���,����c8~`���0����?�|��.)��e`���0��w��?�|���4�����O�|�S?����	�O����X>�i#p�Ы������#���?�|���Q�����O�|��
?����	�O�u���X>�i�1l�r����	�O{����X>�iw7p����'W��l_���٢H��I���ER��%M��&�b�睍G?��7r�iS���O;��~�t���ޝ#��6�9��[���m.G?�O96m�ig̻ήac�3����������p5v�1�:�J�o̿�NNc�[�1�:��o̿�^Cc�󯳿�������3r����4�?��m�hޟ{�~��������������I?hx�ޟ�3���xc�_8�o��g�a��+����p�6ޘ~���j�1�.��7�߅3������p�6ޘ�����=���3G�O���/��^�����@�ߖ��z���}��w4��kMn-��V(��RY��N�0D�P�87klDEr:������'1D !��LH���Cr:�����Ώ1D !�SnHȵ�xP�)����@J��>*�>5���a:T�&>,F&X�X�F)��i��`�[`��ZGb��p�q��k�+�	V�=����\�AL�:�qpX��)8JɵW@L�:�au��ګ  &X��:�Rr����{XG)���Ȏ��x
��(%m�c�]I�]J���V�QJ�N���)�������	V�SXG)i{��XG)i��XG)i��8�8��XG)�R��XG)�t��XG)��i�W?�:���8JI��`u<��q��.E�1���}�	������t"�	V�3XG)�r9���:�R�e]0&X�au�Oi����~p�v�BU(�Bau��*@�*0�V����tu \W�PX]yڵ�
�+�U(��wQ�z���PX�<���^'�0X���(����@�D��*VW�vE����`
�+O���U�qe�
�Օ�]T���2X�ª�s��qQh�C��6sbKr]$���]�1^�q^Z�����r��V8�z�<'�F����ω-ǅQh�C�k8��81
�phu-'�7F���)�Ė��(�¡յ1��r\�V8��Ƈ��ǗQh�C�k�8���2
�phu�'��o�H_�q|���2��eZ���8Nl9��B+Z]�ǉ-ǗQh�C�k9���2
�phum%'�_F����Ė��(�¡յ���r|�V8��f�scǗQh�C�k�9���2
�phu5'�_F����Ėt�"�vE�/K9�,��2
�phum>'�_F����Ė��(�¡�^	��r|�V8���[�/��
�V{Wpb��eZ��jJlǗQh�C��D8���2
�ph�'
'�_F���v�Ė��(�¡�5�ؒV����q|Y�����eZ��j� Nl9��B+Z�}ĉ-ǗQh�C�=�8���2
�ph�'�_F���Ԣ�6��2
�ph�7'�_F���8�Ė��(�¡�^m��r|�V8��s�[�/��
�V{�qbK��Aj���eǗe_F���2�Ė��(�¡՞���r|�V8��[�[�/��
�V{dRb�s|�V8���[�/��
�V{�rb��eZF�e�h_���E�eM���-��.iR_7yHs?���y�JOoڑ*=�dG�������y{�JO��*=ݭG�������Az�JO��YJ^L��m�:V��}[����dp��ce09ܷM�XL�m�9VT�1YܷK�XL��9V��};.���dq߾�_d˅�B��!KB�\2����׳�<s3_I�>��r5��\M�A*W3x�J��y|����#U��-�f�A�j�R����T�&� L�^�G��d��y�0L�^�G��Z���`R��<b�&���#�U=L_�G��d��y�0L_�G��d��y�0L��Omg���MXTb�y��[�r�-�վ��}��;~��4��]�~
8~���kgM"��kg`"��kgs"��kg�"��kg�"��kg�"��kg�"��kg�"��kg�"��;��1%W�qeV�V�QJ�`d0L��-��Rr��a��o�p��;�?���������b�`u���8J�3�	7��M�au���8J��`�`u���8J��X`�`u���8J���`�`u���8J���`�8����:�R�>k0&ܕܥXOau����`L�:���8JI�/��`u<��q�����1��x��q�����1��x��q���3�1ᮉ�.���x��q�����1��x��q���9�1��x��q�����}�������t7�	V�3XG)�a��M�כ�:���8JI�w`u<��q���'�1��x��(%]�c���V���ƯE�uD���T��*VWv�9�U�qe�
�Օ�5�hU`\�Baue��ZW�PX��ĵ�r�PX�<��N�H�Ba�sJ\;�f `�
�Օ�>3hU`\�Baue��ZW�PX]��/�Vƕ�*V�'�c8��B+Z���[��"�.�������
�V�5�Ė�(�¡�{�9��80
�ph��Nl9.�B+Z]���-ǉQh�C�k18��1
�phuM	'�GF�����Ė��(�¡�5>�/8��B+Z]�ĉ-ǗQh�C�k�8�%}#F�J���<Ǘy�/��
�V��qb��eZ���Z>Nl9��B+Z]�ȉ-ǗQh�C�k+9���2
�phu�('�_F���u�Ė��(�¡�5���8��B+Z]{̉-ǗQh�C�k�9���2
�phu-8'���I�+r|Y��e)ǗQh�C�k�9���2
�ph�� '�_F���J�Ė��(�¡՞��r|�V8�ڻ�[�/��
�V{pPb8��B+Z�%-ǗQh�C�=Q8���2
�ph��'�_F�����Ė��������Ǘ�/��
�V{qb��eZ��j�#Nl9��B+Z��ĉ-ǗQh�C���8���2
�ph��%�ǗQh�C���8���2
�ph��'�_F���j�Ė��(�¡՞s��r|�V8��;�[R�R��/�8�,��2
�ph��!'�_F���d�Ė��(�¡�ޒ��r|�V8��#�ۜ��(�¡�^���r|�V8�ڳ�[�/���0�/{E��e~�(�,k�$�n�TupI����C���y�>�#UzzӎT��&;R����H����#Uzze�T��n=R���H���#Uzz>��:P�b��o�ױ2����Zu�&��60+���mB��`��o3α2����]*��`��o/ȱ2�,��qq�&���5�"�X.$�H�Yr�ټ^&���癛�J��y� ��9<H�j
R����T�&� ���;H�j�R����T�&� L�^�G��d��y�0L�^�G��d��y�0L_�G��d��y�0P�d��y�0L_�G��d��y�0L��}[��y��o�_�#���\տL�����j�<���j���jSnwu��ܽ|i8�?������}i��ً���o]{Ě^>�������O�k�n�)Qm�s��2�ƃ�����ן���#K�����n����) �]+|��lˇ}�o��ӿ�������|\Փ����9Li͠��;�e�J�Pb��v(��k/�)���Td�0K��R���,��KUF
��k/u)���Tf�0K��R���,���U̬����fw�XxR�S#���O��PaPb��p5����(�vw�k� TZ�Z��;\�r ��T[��;\��r ��GLW��&�vw��n� �S��vw��o� �S��vw�j����PO�����h�i
��vm#
�@�� @=M�Ԯ���z��]C[8 �4�S����p �i �S���4p �i �S����p ��".��i �S���+p �i �S����p �i �S���W\���PO�ڶ������5����K*@=� �Ԯ�K��z��]C�z8 �4�S��.!p �i��]���~;��qz�u�&=�	�ϕ���8=H��|�segy8N?,���\�iͅӃ��'`��7�����2�_,������No-����	�/������2�_,���\�i��Ӄ��'`>Wv�a�� ���	�ϕ��W8=H��|�ӻ�h�
�P��D��B�6�CmD�D���&�[]�1D�0��	��\tюL(hB��C�+
�P�F��L���&�{��1D�0��	�>tt�L(hB��C�K
�P��G_�F�0��	u�:�h�&4���@���	�+�O�h���>L(hB]!ڧ�	M�ku�1D�0��	u�:�h�&4���B��S���&��]��}
�PЄ�6C�O
�P�աoA�0��	uM :�h�&4��gD��S���&Ե������ޅ�))ڧ�h�&4���E��S���&�����}
�PЄ��C�O
�P�M�c��)`BA�ot�>L(hB]��a@�0��	u�=:�h�&4��	@��S���&���}
�PЄڟC�J�R�O	h��>L(hB틁�!ڧ�	M�==�1D�0��	�	:�h�&4��RA��S���&�>0�fh�&4���A��S���&��;��}
�PЄ�;C�O
�P��c��)`BAj�&t������>%C���S���&�^Y��}
�PЄ��C�O
�P{��c��)`BAj5ps�O
�P{ác��)`BAj_;t�>L(��l����٢H��I���ER��%M��&�b���G���&9��Sp��NoՑ�;=QG���29�Ӄt��N�Б�;=?G�����?��f`w׵���nl6V���ݭ��
X�y�Xk&v��+`���L��,5V���ݽ��
X3��{�Xk&v�+���D4�B���8�B���̣�㾼w�H�	:h���4�Bzo��Kg�a���t�&`��Kg�a��0k^:c�&�3��:e��Kg�a�L�t�&`��Kg�a�L�t�&`����}i/�'@����C�~��|����������!���ˉ�G��4�C����y�=��g�w�Ǵꑢ��+z��Ѣ��/:@t�����^Gx�u��^Gx�:�����:��������a<>�M�׏����Mu&.����Г��a��ty�ϯ���4��xK|Rg	P�Yz�(��9b!�O3k���/����&X7�&�5��A�Cn���S����>��J��T�u��Yn���a���^������2��E��׬L���3(?-��r���?�E?��Q��rڇ~�m��~�h��A��>����&�i��Y�/�݆0}��g�^ �ʚ��1���2�,�7ŲH�i���i��"��U��g��/��})���"��6��РR;��VQ�:�N����v�us|�/%�/��t��E^߾�t�B߆��������{�\�s���E87;\�ʉK�����-����U�?,��5gn*G��0m+��k��K[����j�睶j�G��׾ј$���ķ=,=PfQ落Ӟ�iR��nvL�����Y!ӣb���i�eꏉ=��>ܘ=�<?>�o3	/2��_8��V���y̥����Qfv�0�2S�ݧ9wTq��gG���Q�Vʋd�^1W�L�OI��=*�>����ai�N�/)��c�It������Z�4��s��=Js��0�cj����1���?˟JY�\P9���1����>1q���~�sq{ݖ����?����s��ȋ��3�w��~�hE�G>�w��O��m���o}�v�s�~����R��=nV��1�{x�}����;�[V�&>�����zX�����v��W�&��}<�Ī���<.���q��.<=�	ɮ~\m� ��'�$�g/���5�ODHe��#O�?>��Ypi2�2�L��6���9L�f���������u���ڒj���b�7���̈pH�3CϤų�C�w\�7�v���'/��R�i���}#��ȟ��ۘ#��R��N{����tk�Ȟ��������y�6ʮgD��i߈,�yb�z�����OOğ۞'������oD�{��a�_�	o��)˧���nv�^����������~������dU���"�tZ%�G�w�&�|���vA�l�K���r���
�����7Ǳ�bܴ�e�j��t�̦�L�ʅ�By<��c����+�����"��8��L��N\.E��y�|��<������`��*�"�R%3/!N��P̧�P���|�f�ߍJ|c��S���N�~�Z�O��*��,�}�ǟ�Y���]����4�"�f�B�u��m���7�'*��^�&m�:N=��YN�y�('�4��2�dQ�gT�^o��4�Z�U����i
�1�R$U���,�Ki����W���qz>��U�s��m����V���]����q�m?=�OYr<��������v��}]������6{O�1���r�n��ڋ���?*���it5�:9,���W������F�SߗoE�ϋڻ8Zd:V��,M�.�Y�5ӐW��΢��*��V_��d�U,1�4��e����[�X�󪈧�,���Y��X�$��l>[�E?����8������yh���_���ëW������&��������̍}��5�7����qs��'����ݪZ��7?�6_�������>�h_`�ݞ�[�6g�w�}S�z��ً��I�~���իW�?5�����8�ۯ��o�P��77u�������!?6�f����o���P��K/}�Й����sG�6���
��M��#��{��G��Z�e��I�*��w�z�F��˃o��Oo��4�2��ӡ���U�j�������f���U�����A/o|����f�o�S�!I��k��a�9��r��fS�Q{a���U�~�J�<<Γ��`�/�ġ�oc��P�ߴZ45������۩��>z�R�0��~�i�4���3G�g'�/G���V���c,�1���J�DۀSEp���RE�����T	~H�<?ʻ������Y<l`��&P�����q��:V���;9h�aG�˧+�Ǐ.;_N����<x>�z�s�՟.i�T���~��K_�Ń��;6]��.Ϗ�şσg��֗.:�Z���/���B���1�������V��j����o��[5/_�|�?PK   g�X8�w���  ��  /   images/219287a5-9258-450b-9fa3-793f4dcddf2e.pngt�eT]ݒ6�qww���=����7���N$xpw���!���s�����������%O�ڟ�eP	A ����*�A���#���'@��,��)F��A\R&�	ܥ��՜,ݽL\-@^^^,6�vnf&�,N�V'�� 9HNRL�;�軗7��@G��#WX���&$2RU=
�(�h�OLR���
	B�X�*�>�z�hP��2���H���;�G/��Ga�������0UD#�� �|y)_k%�E�	n!|�Q�xH��:o�'
�󊳡k���AV��Ehl�atܽ�V�}�-£�z��4*�����R��[C��sN,�4����t�P��P1�s��k�a��[��9Uӳ��$ceoZ���Hd��nD�N���z]`bX��;��n>��v���*/2��Ю+D�Ѕf2g��
ZU#��*�*�Ɏ�$�r\�gq+�R]�P��blz��r"�V�m�BO���N�J�Ӕ1>��Ptǟ��.�;���r84(#!*&S�����C�,�g�"��oá�l�mI�b��k�}�*[�:���rF�չ&�!O1ogX���@*�n��^i���KtW�U�,�p��d��v+�)tpʊ��мb�!�2�L��uh<�V?y�M P��<�	���?Sby�J������Hb��<խ:9�c��Qv|З�͉�c
�:���9�	�(���)HBOT�����p-��b��A�Aa���b��HȣqH�_�ۃ�#J��s�'��L�	B�r6���ul4{��x��i����=8�O�\QF	A�|�&�
>�9�Kv�mb�U��tbDev;ORq�`�o�Y����v�G�P��ˡ���h�3irq2��[�&�����l ��E�lP�骟Mߑ�J��2��E���b�RE��/��m�*�t�jz�Ƞ�*�M�'.a�+F0�6@��.g,S�P�xZ ^rߍ�!*���,�)e�q}	�z�"y�L�bTtE�Bs��$g.������u⾂)c���.ȉ@�F���t�>�b�XC��433�024rQ�I��ʑ��������H���L8�X�o\�8�qgt�w�t��|h7��*�� 	�O���bcP�����?y$S�>���Gb�gT2R��dܕ�u��|F�S`��Gz��)K�jY^��2��Fl������\���o\��8�\G�!�1&h�A�����m�"5��#��
�A��x���+n�<X~&Aڷ�cQ���V!'�졅��rx��}�Elv�4{↽) ����o+~i��K�#\�o�XF#��`�kL����0�TO-�;����"�Ck�������G�f����`b/ ��M��vgC�1|���Ou+�����ܕ�+nR�Q�1�.��7 f ��̫Č_��zE�E7�bc��v�ɑ�*�j	n�g�_&8s�S�J\Y`4`��J����g5%e����5�
D�6'9�eS!�G0���s��s�~�ԗd*@���%	� �[��J���0��)�nV���ݪ4UY$���G��6)���Tư�:�&�X?Ƌ�j����^�bs�7ߺ
J�M�i�S�ZV�:h�+zO�8�֕e�8DlF0�}G�SM.=4)r�1Mw�7��S2��Hb��)UG��>b#
��+0�B��6ϸ�������Y���Q�I��F�b�O��&�Y#
忶�&�A4Պ�@퉲��%�̇���5(b���(����7_�,�r��w[|�6�.$��W["3-��������'27DMbɥGg"yS�&�A(�3`qe�Qѩ�,?��ol
�Mb�KN�P�B��L�V���]Y �@�q"׬���p� �Lg�6gn�::$���/n�(��SʒĴ42��FE}VXD) QJ�|� �7�J&tQ��F>m�wzȥgg"��$�C�5	�:4iF��6/�$r��H{��3p�H�M���T���n^���ռ3 ��'C�h��GT�`�i��m�C
F7�;�V�~_f���BV�?�䪜B9����[�Ҝ������B�t���a܅�oV�ҷqi�t���a؅�%۬��/Z�-����:�B��/�֨�`q�{`9���@��"�k꿚��]�w�����C��0����$F��}�I����·�T��Qs�6M�C1��sX�n��V ��M��Bz�5���&�"\�/}Oto��#�ŋo�x4�3SHI��oWC=�/��@p�r�5�4�{f:�Yᖧ�d"�r4+���({I� | �B �!�{8��;�>��X�@;��Z,��l�qp�.����+����VR&���T�vL�Ц�ۅ���N�<��ٗOt^|g@������s�<�
�K�\�*���VT&�̿��,�F�ㆹ�-�P��4���:��Hy��e�=��f��Y���Vκ�f[j�!�Y<�&�}�R��u�r������V�v�Rݩ�����Ue�Yeu �d�R�{g`���y.�ddd��H��=�s����=q8���^�"l,��R���FJ�@?m��a\��-a*��T*ӛոe�:���:�
p�Z��A�f��T�]Hj�b���T@��1 �ah�i�d"�������3��h����_�|x���o��D�_�Ə��*>KR��뱖CJ�$2��v��fX�4�S}�Q:Q��:pEsR�#c\M�5�2k�̰�CK���������m|+'�dQ���^�(�r";E����;:���E�8j{�4Qsz $M�G�j�@�ä9�ˬ�Y	�׵�w��z�׾���>��h���;�Y'�(ݕ�Q�1gJ���,7f�O��g<C.��$d�� OǋG������Rl���f\m)ts�F��O���s��֥8=�҆�w6 ���]s�6���>�<|h�^��>�R�7.`(��a���gf\�����Rl"�V�D�J��Qh�1�<��֊̰Je��8��1�f��<�mUEH�'W�]er�X�A��hv���N��B9��vWC��i���N�12�X*�f�J���.�����ԩ+��N�cN+��KG#î�t���%��5T�����?�t�$CW�n	(��-�z�L�OѼ.��ƕ1�������(�Q^(}��v��I���(/�-c- 9�?y�]��ha?�R���+3����'�>ﰸ���d���z�a����^=�,�k� AP �W,��:O�7dcrP��8.^j�9>2lh�1�/	x����V
ퟛM�J�����.}񈌓�A"� �0Ɂ�^��U�3z���s������
�7���L������.CF���*�Ġ�Vc�儬vݔsZ��R$�2����`��3� g�)��� 敜�[�����^�3�<AL�J��r�ވG�G�>Ձ�ߴ���l)O�mJҷ,��v� >�z.Fe[$o�s<�F�,�xL��̾����}}��6�q	5����%��1��ŵ�4���=�HB��^%�m�������ԫ��~��ch5�՛�%��YCY펈��X���]�łM�&�"$�,��?�E��.����)��V���4R�\�nӱ�N���l��Nz�h77DȚ�����>9ѫ��߹���F��|�Q���ex!��z*�=
$��_� �y�tʹ�ǈ�Q�L	y�T�sNi�9��Ґ� �yM�7��)O;���)�̲�߽(&'�������W��;f�����=�`A�ivj�=KAͻ5����t���-P�G�:d�f`,��y��Wߞ�U l�x�;Eؗ��`c��(�q�ÕL������Cp5�7��q�E���4�e��F�R��P7�ݚ!U�h�Zz�c�����\���c��?v�cm|��������b^�_�zG��_���5泩�][5��q�J�.VVˣ��A��Q�~F���5��������+�,y/�N;�C1�XSLf/&�&�}��E���V��`��ow6wn��vj��ߚ̳ 8���[O���lԼ_F�%m�[y�U\��K/�u��FXAξ�S�^��xA��F��;��Ki�M�[U��۸#��j�$�mE=ul���Ҏjg�2hɶ�cA�%��eO���ǒg ��Ӂg�����U��մ�*�^U,�3g�{i��b�[����CvR3)��,��r{��i�S��'2�'�Q���R�>��j߻]��
���9((�=7�g�'�¾�V���BJ`^���#�J	-$Xy���	8S�wM��d�0��z�K��}�d+S��}xd�&��mH���@�0.�6�-ǭ��5�1G-,g@��s�boF��g��.����*D��+�A��P:�a�״f.��f���i0�!����J4�BM����JZ��)��?Ի� >f1ev���؜	R��؅l'=JD�6�lFnT��`�oщv#Y"#em�>���ə�*�
��UM_�_�2�pSC�Sx0��*68�]54_��� ��T�V����V���:�>���&L_�Ru��0�,�Ϩb����k�Բ�u�w-���X���Q���l�?T��S�bQ1#.�u�m���@�T����|�9��7v�ޣ2�P	���_X�/�R�j"�O��Q�����A�k�	)i�gR���]
�%?L�{��g���v�x����ZT�!5�%+��ɿ8�Z�~��"E�UW��$ ��+ʊ1�tw�X '�A�=�b�B�Uٌ���xl.a������|0	���	��G/S"kCax@��8�*�c���C|��	�z��7�7����� .�M����׽/w.�}�$���U�y)��>��US�PV�js��qe�dy��yo��<���L��F��E��|Yj<Z�b�z���0o*��O�Ƀ�4P;�v)�֒r��FTIw��y#�s2�6�N���"c��]ψy#ɟ���b���٢/"�l���۸����IS�0����a:?��B&)bl�M�<��pT?G=)Z���#����Ŷ��4ۍ�l;tXW~L�/7��볝�ϩ��t��_�"c; �������«�_~�_#�k��&+���>Be+�o�!mX�rX���x��hޔu)���2�B��H�ĭ�g�uë����j`��R�X+m��צ[�ւVǫ��:<�p���gtU_�(䋎��pP����}nMIj��?��L�A��n�?85�2�?�#��WQ1:��C&1�28j$�{tx�%&��\�8fvW�<�)$�S����:������?��S�h��#mx%�s���W��9�K�w�j���m�*�� J2R��vx!��!]���#敗�緵�Ƿ�����}W��o�!�#�x��/$�eX�-{H"�UܯAJh���<��hEq��;��OA~�]��0��ĢB'$9��j1��h}d��8���3���šg�:�c��W��[�A�$����}��]�����d��_?��"�o��O�y[�C�0�������Q���+�^ppMu`��7� hH��������������+����J�ץ!����M��'��H��S��?Kϐǻ���gI�1�kՋ���B�b�u�8�4R݈q����#HM75��Z���M7w��F�5���͌Q��^r��׫	�m�v�i���93�Ot���_��.��ٟ��.����8W��[�ǘ��(W�Df
��R�Ո�gL"C��v+�Iv���Ý�x"�{H;��l��9����R���`��ߩ�N��y|o^��ؓ�EҪ:�+�#��ɶ�
��*�K��Q;��8�1x��YU��B^¹���yR�a�BA��/o9��MqxW���>�@}:T	E��M��n�&��V:���g�_l�|0Q��m*�n�&���2���mSeR�&�cx�z����	���6�Tx�S��i��=���?������O
�bc��0�\8���L�"�ˋ�n3���t�O�,H�e�H@~W}͏��P��V�+�T`xr)�TOLb����T\���1 HWQ��ʃ}��ԫ�ŝx�1����y?|'x��.���٨�+�P���z1.�����>*L�,쯅�$~��"]O��N$���p��u����"NF5{�Q�m�O������MI����j�d>�u$9��|g� �h	�}����,-�\m���\ѦqV���M����/���7n'J)��Ts�w!�S�5��aE���\Yr��*�<�'O11�Pc&��ߜ�
K����Ǝ~��NB������Q�����@uf[߿�W.�`���Z�⤀�L$:����m��O���|o��{Ԣ�""8ȃi�M���á���wm������c����䚩��;�tr�e�Į��T�q���6I'� �4�u����2 W�rY rSin�����_9E0���4J���	v�'\5��N�ˠ�*�3(�� �Tߵq7F����B�'^-��3��������ej��RSv� ��>���o�M#1���|#.xmon��0=�3F��:�PE&��^BM~�������T7�&�fWr/9/�1�m������e�`YK� �.�k���0��]�+�#0a��V2�ZBh����#�cO��U���#!N�`¨�Tu������]Sܽ��K]Y��#�7�?N$��?����W�IT&Ҡ��63�j�yn)���$}�><熶u�ߚ���T��.���;7!U�
c90\��mx�.IM-�g��k1��w�v��7e�[��TL:�����!�+:��i3���8`�f��M&�VH 3�[�d��$}̯�"�, ��#w�ϔ�?�bcqo�)�QL�6�2��3���jԂ?�vk�i֦��ja�IM��qb������(�$P�N���Ŧ�J�w��M5�-p����?�Wd�C�o*����ȝ%��3�TjJ��f|5�m��,�T�w+X|x� W7���*�C����N.�8
T4��}�T��	����6�+yg����f�z��T�/���*F-zj��&sU��/��3I,/��)v!�|�ĺ�t�=�47�bj����k��4wv�H[9<�1�ރm/<�R`���T`S��c����b�3�����L��4�	5-��D��� �e�w+z=��	�N%!���N����j��%�r��O>N���8?�)��I,?3�d����K��j��J#�<4�b�h���L~��S
��\��v��
-/<=`4��i��7<l�*ڨ"R�,�r�UFU���n#Ü���k��;�D<��A�����j��} e\@��Ж�R�����Sh�lzU ��t�jv�ۓS&'�V���d.�	0��ߋ�o���}�H�c��ešA���i�U�����C?O'�ԑ�Lp������r+�P��5b3��g��zz���5~b���`���q���I9q�}
l��J0�L�r]E�1�c��᪓��?�=��o�OzU��s£�NG�v1\D"6E:���a�^X����D5hU��W��L��s�DV`�0�r��-p�g1�H{�@��]t���T�� 2U����5(gd@����K�*iL\}G�"����pQ�2l��+}&�Z���9lݠ���ʑD�|�Uҁ��[bed��Q��Y{ű<O �FU�:��	�?���c?��T��*�h�,I�@$7�'�eɪ�$�XL5H�����2	h�8��?n����o���Lf(�o��0�i�8�pK�^�����ȑ��sa$�B�;�?s�*A⃗�,����ݓV@څ[�(�!��wJ��|ğ����3���o�6Y�e��&���cp}��~�#����?ҵ�"�&�*��fETО}��tխ�Dq�Se!=��M2[ĉ�����k��]��y��64�Y뱱�p����������3��A��f&�\�$J�YOW_]��#��ʏ�t�)�s��3}�-��eHM�]�?�-��fkOn�M�J09���J�i9*���Y%�"��䵂ڙ�w��@wf�A|��x����j�H�rn�j[*�q�l���#jzS�B_��U���T,w��`�OM�ٻN��pC�C���	I:�*�,b���:Y� �C��<��PQV�=a��|'�<�B��.e�����a%�i��2w��]o���>�{�S��u�3�1�Nc���){��把g7�p���̑�	�B������Kc�����2�ʵ��v��[��'vz�#Ó���}8DÚ�k�z�1�ᰐ����Yko#nc��L���I���%�����h�v�B,5X���%���T:Ɗ���H�u�����p������!��r%H��c}�x`s�h|���ߓ��\*ɰ���Jl+��c�@
�|�z��f���-�&��]�i[L�!���`	���q�yrb��㘰�Q�C::����r���l*�!%geЧ5�f��O�=�;�mC�ެ����S_M�J2�����(�k�#�Ō���t�3�%��e�WG��
<�W��_U�s������c�k�.�)��'m���n`0��U���i`���/Nmp{?��g��no�t��\� Ǩ�F0����x�B8�O�B7;!&Nx3���1��
��>�U7�R�K�����R5��w��~>�%_��`�G���(z�m/-��pC@%��ij�H����$�E��OFH4Xj�J���A$���k~$�e�}&|3.�G��ʺ5?d_�{��z� �<����z$�\-�si)s�`v6_C�p���]^-8��h��yzv��{�[e��aq}���:�wvgW��m~�?l�do���ZN�]�ϝ/}�x�����ڵdM�m%�H:�7ܵq)h�MVk�>�{��t꽼�\"s.(%WLjU�j�֥VW�e@�K�9ޙ}��'�	f�|���-����͍���(�Z�s(�r�ӼA�D�����56v��9Ͻ�YMڈ�-@h��=�(K��$|!����]ܗ�ά����n&Ґ�`�I��~R��I3�ý�j�'^N��,��E���ƞ�I(����	"��� ??�����v8	-81�/�̎M�sj�,p�.���d���O��亜�D8f�����fM� O,�� �GAUϓ���4�2�0:���b�`�q��]O���]�Y��`� �E8�{��S��Yy5��l��e�)Q�I�։���3��+�b�{�����3��fx`lltY/�A���������zW�w~�Y=hn:��፛?�b~d<��:��S��u3U�m�U��G���������A��h�� +�~��*�F��4 ����J5'!������ta������yn�
e
�0��62�W?t�oQ.ѱV@Vn,?*+�c	�s��T)i	�����"P �{�-ݜ�c5e��F��{Z��mﻡ���
���ۀ L;L:O���}b���oa���{j�ߝ� ����dtB���eѼn7��pM�5�����{���Hd���l(��`�A��LBQMD�F|�iw���i��-�b]��͂��p��P�nY@���cT_�.Ywo�������jID�bh�y�Q((��}����h���}��� !Gۈ@�ȁV���C�p�0πɽմ��j��{�[�Ht�m4oJ lŘ�Ǽ�T�?�*^[de%y>ɐdS;&�'M�����t �W/ט~R�~�k��%�؛̓BDT�l{U�<�[��%�����i_ߩl
��B��E����zi8=kY�v��$�K���|ۙ#2���dɳ��i����@���;��� [L3À
��&��ۆt��5%�e����c�~ N<T�9y�Vo=+X��Ei���g#���\�d�9��Čp3�ݦp}e�3��>}Zy�N��z2f�m�c�~��aF�>KȌ��;�Κ�̘ؼ����c`H�ҙ8d��	������e����x�#�l�C`6�Ҟ���mWge���Z�CPu>ts���R�%��Ȧc��]�W��==��k��0X[=׮ߓ��N�|��+�^b ���o�Z_G)�3W��j�92�l{(詭��y:����n<���&{M��acpxHBE� �P*�&�����gO����q�%9D�Σ��
^:�1���,e?���LwCM][��iwD�v1<r53�$u>��BU�ҿ��_'�$\�R5�9�v5�7;}w;�m {���[���G{��nD��-���l�^6�:nj��ã��7�=��[�݈��ib�IERCٱJO�&�۩�.�4�-H&?��7RK�-����w�Ԓ�c�����(B��̯"��
�������Aۙ�0��먝���gdЊo�	�˪��U����z�·����c� �_\�k���c�-�2VpC��e
zo0�����1Ds����s^��Og:��f�h/�[��xU6���#���޼��ɞD�-'/H�\��a�l���}I� �G&�j�t�sK��g�bW��\#�=�� ei�΍��4���� Ʋ����VI(����u�f.	����I�����k}���ʅ��-�v�:��I�Ѯ����<����x�=�鰘#�����l���6�js���T�i�N"��W{��j�h��+�ox��̻ C���)ѓs�E�pzx�͝]��q��J��͙��{j�a���j��+��l"��΄.��+�[��9��s�*����P���]��z�s���fu�t��'�ZY�5��/4m>��$�.ӎ��`���{'�ǋY~V�R؛�(��O&}��g����N���ڐ/6�v=f��(9Tl�rXQ��� }B>�9�6b�sd@%��� B���y2W=�.^�^Þb&�^ԫ���Y��ؗ"�h�ܪf7�I����d��l֕��t���?�3��8S�����Y�󭆊��x�^pNJ����1��Yǂ���1�:s~�������@�����h�a�b��%�zh�a2��hOzfl���G�e��ӟ�e&�58��Z� R%v����-���$�O�_T��s�M�e�>�{���{��Q�7��h�9 �>..*✕=�[j&d�7bz\x��P��r$�Y������Ck�7ڌ��>uK��d��|�6�ǯ���������q��L����9Z����q�j[��6�.BZ6�_��\�� 0�콳6�������;�|�J������}y̞ޜ���ޟ����t
����Vj��'a�׈�BW����=�@|k9�4�W�G�,q��n��~ӺM@���~}v�EY�΁@�U����B��ŭ�AY��―��=�Ps}��V�m�E�3�����H@�����S~~˄�4��|u�խ��-�����Q7�L�fTE\�|9������� �*˻N�@�)��
�|�+˔��x���P�M���\��������6Na;���ĵ@$b���d��q�7n}��1�^���cBW�y�=�_�^絶����*���q������� ��ǣ�]x�� �҉��Z�>kN����2V��%z��d�t�󅹌���Y�ـd��<؍//�Z���A���v;�>-fUy���yz+��ܾo��sK3*���/�&Z<6�S4:�s�U�V;�����<�J(&MF�'_��n�&׋�ʭ@��?i6�������nk 2�֤�b3�>��
\P�\�=~������>�DG;X���O{E>_ �
�UV��@j�m�A�����p7-�������GY�q��^
���?�n/�\Q��Y���ڒ���|i�"C����/� k�C�6" 
���9�N򕡕	�8��IZ�x�iO��G��0gD���
@ț��޷@����^h����B�o���v����S&����!h�]�" �4i ,[ϐ�����{Y�qc�&[BA�2X��8�x{�!<H�'�zά�G
 4�;�r����� 5ҷϘ�4��j<y$�ueB�w��P�ԍ�p!&���ߓ�<Jb��^��R�ޏ'l��P��h�-'-�)�8]M �L4���ͬ
��?u�b+��q���o�̑-nAy�K#5S�a,�ˁD���鱃7Y��[�=��Lޯ��ָ��h���L����ۑ&q�}�[݄ɞ�Qvv<T��n^��&JF|�r����H�����Wr�;�h|��"}EH"r&�0H4�L~\����
��.�E,��v�_<��9�B�Q�8����J_~%�P�n�h��l��e�����gN�,ը�
�����.��w�����5&s~��P�P1{�7^�D�v�����P)����C$�������:R�6z5$<��!�~$�����h���[S��y���Upm�JI\��k�6�f��A�Ɵ���vF<�?��;�q7L�]�M�1��b�R������ŝk��V3���WR/旘��Ɍ`�jQ��J:�t�$A��[�8�=��<����Dc�z4:���O�P���t�/�>�.�ߜJ�ޕ�:��1�d
�i�a�,�����3�7�8jH{�,��.��=�v�GY�-{�ޏ���~n��5��ΠMN �4��z1=o���m�ZG�.�l�An�[������`�!v��� t�0P޶y������{|;n�
v�E~#�����-���4��[�?IO\�X��t��S�����\p��oHa�t5�b-Էd�u��U�:"�4�>�t0'�Glǭp����<���r-�چ�p4}�<a!��a�|yFu|��K��N��z�  ��n����>:Z�ĥ���b�M9����BL�\�������#�~ �i]���]8�ݏ�:r{��y�eN`f3{#ާ+���k!����U&�Lа}Z·:�5?Q0HqÞ#ޗ�o!�]FU��8�5��w�TqKq_}�	c	I�|R�D��&��_�l৕/���Om��w;d��0�wfKb�����y�(�(u��\��u���Fa�������L�A�\�_��jP�bPihX����k�!��I�y�eA�9�f[j�3%�_����M�T?u�>��ru���c}/:Bz��Q��υ3��=�4�d�g��0&��?�>m���FȌ2[b���6��6`���(����^8��#���l������۬��&__d�s��_��ӎ�٘*���oI��8M��,����i$�5#�#�� �c��,��|A����2Oӟ�&�'�6��,s���z�����/;�G���.�Y-d�}VHYݍ�Pg�Id+q�Q
�}���3��J2��F:弜�z;�yVU��������.g>�u���@�;r���L����,�ɣ�DԏM�Z;��F��J�IXb���cS��ɍ7�*�RX������+�X��Y�_��a����������|xg��q�7�u�c�~C�eY����C
�]@҄7��p�5�4���]}��lɑ��
yv�\GG?��fz~��*�Ts��x�
���u�]�k�W��Fч�	�Q�������W��׷h+��M�hftK�3<���S����7��|!��~�y����bIc� �v�w��cb�����S�J������Q�������X�Сň��XI��퇇$�߼H���~� P(u��q�������T�L����9�dm�ë|fUr:Q�QX+d�^d$���B����QX)�q�G�+rrr�J��x��u/�}[��!iD���[���KQmt"�Xͣ|��5��]���~�^nc�u��l��c0J�o<�C�����E�k~	�o0嚱{E�>�L�Dp*:j0��_LE>�Fq�o�S��fKگV��ގ��yk����銀޷d,' ���!�
m�37�^�4�1��8;��]rfd�:̌X2�bo	u�H����E�C ����&�2�2�W�uE�J]��\i)I�av�|=#�Z���ݬF���1��Vxh8��{�l������ޘ���������p�����f��_�l�� ���znl���A��C�2&�V���7+��!����f���9\��M{����-����>D�"��[=Ku�@5�i�H���7�8L����:�۶0���/.��3:���fޓ�T�D��b�e��[���~\��S����%@�����͔!"����G%����$z�)bw&�v��'ۆ��7�i	�M�T���"����c��jD������LF�F��
�!�4�[t���͐�wFd�o�T6��s���~���f�Q�I�s�����M�
L	i�G�Gٿ�T��'��ʴ��~r��ƟLw\�)����\uN�@���G���M�s���	�̥�M������[M	]\Y��U��d�2�a��$qv�� �<ǁݑ��
hV�o��(H#^X�@T�d��kl��ZW\G���\�D���Q�>6
Ѣe|ǈ�R|Ȃiߓ�_�Y]>�h/��I.��ՙ>�p�g%�-�5 ����g_���&Uӿ�4�(�zs�A؄���ɉ�Vpj�E1���x3�p%1����鈯��vBʅ��F&U(\w��|6a��IhDI|��[�1Z��D��i��q��}]��ߝ,�T�y���ݾy�*�7�*��n�F@�������<���ε�*�22��$~��T��h�s�&]E�Vo(������{}��
��o_H��.O�] k����DhF?�n�YRq8�(vn����0?����`��ƅ�"o�̥��cx���E�Z]���l����@.dd�)M�c���D�L�k/�\�>"Qa��K?6|��q����ff�i�y��XC���Ijq���>�Sg~��hr����ř�N�f٫	ܛ�ݲ��~�1�#��p$�yؾȵ�s�����d5q�=�,���t���iyN��Nj��tL�/�ﶵ���ɉ�e'�����vn�,�·�_Y��s|���~���t���{n0�c�����ŢR:����݂w<L��*�i��\��t~'�>Y��f�aPꔴ^*Uk!��|4�����@�v��A?G
h �����ͣ51���/x�3�I��h�_����7�*V+t��]����F�v�:OLM�}e�$�����Fv.�͒�O�R�<���u�F��㖩��?���h�6.��"���vkR��5�JYhh�5E�W�6Z^���[��)�	�_~���3CB=��9�(5���������� ]<g���������v��8U˕�Ӵ��{�nӺ��o}���
�o5��a���� 2�]�E���5P��cl�n���S�6_!V�}�#��bi�j�h��Vԋ�Qo��8�0㓲��._n���7��aD����C��1���ɱfM7n��k��;].j�k���#2 4q��7ȃ�̝2gM���%�G}3o�C&³j���b����I�Jb�MkZ�i ~ g�>e(�����������ҙ�7/C�Yd�~Z(5�7Ii醆D�*�A����]��X%9�E�Q���w�[�q�WST�A%+�-��/t�b��I��������^�8��X���L�{���EX����`�>�1Y��$���? 8�M��gP�����{�#���"/h���NYn����7�W�$hu�z�KN�B��N��� Ѐ��,l���f�b����gkV��5ӟ4���O�pG��ø��s#�����>����.w|��Q�LBR7:���O�Mݽ)]o������k���s"�ΰ|1:��f2O^�����H4u�zGN_���p�����Z�^�?�x�b��������v��`�<�h]$�89��o����sf�
��2|�S�zE�����e$/p���`��g	�s�0R�ĳ�{q��Ӡ���,NA�����ޯ֓e.uǹ��*����{���_K���qG	�2���eT#��|��Q��N� �3��C�Ņ����[S���hi*��8��L�
e��R���T����sV��3����j�$m�`g�Veۺ��v�R?�<����C[�5x%���`ۊ�pq���"ph����in�/'�t����{0>�����AZ�V���L� d+�4eO��lԨ#��^"��܏�ZK�7�G4�����.5x�Ά5��b}ꁋE��`ShQgͨ���-j�&��v�`VC�+���J��z��9���"�� h��F��Ӷ��D)亢�3�q�$<݀�5D�x!"w
>��+�.�H;�h��/�����{oCۺ-U�縯�q]XX��Rk ����k�ފ�������D �`���.�x����m�%��x	��>�["���y�ǲ��LW*�I4���I��!��)f�� ��G�m@ze	��(ح)��tX��n�cNy��Ǎ4]�?��sH��E �#V��t�Jr��z�/b	b��c�B��;��w���$s=�~s��*U��Sc�����!i�5�����2�;���^.ߏP�Nz�yE��ゞ��=[�9$��y+�y>}7,�mw@^ͼg�����~{����������>xT�ݺ��#15��1�߃K$cv�"�q��O���zn�~�������v�/b}�3H{��]�N%�{5�}������4'ec�L�H+�8�����!u*���)��_�NM6[`!-c�FW_ 
>wH�n>��Xƴ�j��3A&<��CI�G����7 
��D�+:��~�p� �=���,���={��[����0�%N�|���Jj�O< �I�\'V<r��(�p�z���&~��S�e��N���*�xo�*�ǉ�wg5� {�ۏ�'�|�d�.�sc�q�Ƿl�����j���EAT�D���R�w��+H�5� *ED@A@z�%�BT��tBh��Jh���A�s�c�W�=��R�^k�������=�,��jG�Sen��S �ۻ,�K��3�N��|N�!|,�|$�ΜcB�褎wI�7�i�$E/(	��q���������U/����l��mM�˕i���r�)�H!����]ߡ,�-R�P�{�{��{��k�ec�d�4:���Z�~��?����G� �0�Re���d�
߬�SE�#��G��L�X�W��3y��Nڒ^�P&؞y��/D�L]W��ȣn�>H֦���aF񎩯/qB�	h�:�?K���U�O�g���.�nkH�����³�;*�2�3��a�!��G�`8e�5�)�-��q�������u#
��I��`�y�:����t�)Q!��S��N���k�5Ғ=Y]%>r�F����=�q�\��l��h Z����% ��@�I�]���!����	��"���!�6�@ڵ��@w���7�_�C:�M�&��-KFPf�1��!�n� =�A�ۋ�ҋ��Wyy��ӛ�p����5��I��8 ����!�D�����[Op������\���S��P��@���k_zE��I�n~�1]��lI*L~� ���R������BZ�x���p��>v�&�����ʒ���R��K��-�~�D�b�� '�<9��?��E��:'�o�����}��H�N�C�>}{J�F�iL��9��  p�Z�G���^m�J6�ӏ�e����؊�zb�4_�2������G*�.s�����}��0إ@�$��;����*ʎ<&d�g����[Q �lK��'^b�Wb�h�n0]�<�����e4���O{�:�^���I�J��5X�M@�GV��}��G��c����Z�����ѝ�N��BZ����B�	�|�R(q+z+��F+}ނ�M�jaQ�d��U�|^��g?���6��z��Y���מ�M��<�� 1h[��xu����e`����)BH�$��٘F�r1n���)/�=�qu%XC�+^2߭�R��v3K�1Cu>�=��J;Mͻ��Q����ܹ=��)Q�\�!v���SE�ξ#�gs����R�T�k��}-�i�3_�n7��)T��B�2���=N�뒼���Pza]v�m��ۛx%������/�o_�Rpd��X�ʞs{��@B��ok���N�:�J�}����Cx&�|��5J�qN�) 4�P�W�����[@��(�>WD(jd��.�)t$���Y��T��3�)%|��b������
�>MFq�=U�>~wŤ���1�\AZ(B���_�O
��x����ܰ�i�WPT��n�s�ܴ��#n�Q����!�n��۩xܔ�%�gT��Ǘ��s���H-ҫ�Tgʲ>.O����Q�a���VC=x�{�T�5�jc\��ٍ��X�-
��-[N�6x�ΕbeHvs����A��8-���	e�k����f	����\cD���P�*�:�=.fT�޺k!m�
�F��-l}�W��~��	���Y��#[�ߏ<b���ŉ/	�Emmԛ��&���ў��eԨ|��)�r�_�A��b�a�-RSkH(�	�GB�cas1�A;���U~�0���utr?�\^lK'�`C��wi�\�&���{�dAc��*S?�9����f�w��,J����^>:��,l!�8yC��<w=������))3zњ��:�l�s��:0��ycm��cB�5|����<���7k���b�ל؂�.RK}�?}�]V�����kr�����9��}���d�TT0\��x5�k�g��c2I�ӽۋKK��gU?������\Ն������*�Ŏ^��r$�zq
7vt�UyoF#�RR�wM����I����{��A�C���h��a�J�[��":e�����=8���T���?8��2%���������'r�ˋf�BZ3��BZY�h}�|
��&8�>S�.�o�ͻ���O��'������m}5�c�;X3���m�zb��9J��2R��o�����|% d�xq���_^��y������{��^�'ĿxBxI�⛇2���H�L/>���#y�����jh�~���%�z�i��$�j+�'�פi��c����N�io2j��yCM�y�)&A��|�U���U�~RH�cF�����=$U��A�����$	�����!�ǏWu5�_D�{��F��Ab�8�t����1�1�]�������s�2N����J&�B����'��4-e�*~~�וh4dF�k8SV�֖.oe��~$���v$T��O�/�R��뵠��gМ�:t�JE�Kŏ�c=�&E��i�LaZJJ�������~~Mj�"Y�)Bʱk#%�D$�?+���PX	"I���O��L���&��&�˙6V���1�k���_RR������������G?����=9�cb���ϰ�������y`���ڴL�~�q���}��Xf\mԸ�Sk�����  ���`z積1�=i��^��,,}�Si\�OĬ%RhR�t0�������w$���6J��PEͧ����'����V������X�ii���҇z�'��nP\����*�����3�����Cf�����9�S����k�����;݂�P-���4��O�'8R���Ƿtgc��ua~s�zo�^�ώ���djr%���au�gm�O�jZx`�^�˼����^��n�TD%Eȱp����g��(ی	+/���܄�h�m}��<�J�K����0�d�{L^vo��|؃�6d6�F��ϣ�����N=��ᾒ�;�F�$'����*�ǹ�a�G�5*
� �&�^i�Y���;9�>����4� �t������U	�G���/J��P���b�?��΍'�^�lPT���xM'{�?�ka����%�{.S�'[E��Z��ۛ�cy+L��ʵ�2��y�Q��ڇI�ݶzm���B��Q�Mo�X��՞�Rl����%竤b��;����0�%���	���;�̝�Ȗ~�e&���/���L|�^h'��ш�q�y�3|�1�  iX�z��\; L1 �e�̩ķ���71��qx��C&��_�,��wML����'���k?��ܨ�zb��J�C�p�C�|��#��>�8o�l�d��P�YF��wMsҞ=��h4!є�bY��棯�^X2�'m���a��dK�n�NJկO��t��ĝ�QKL��t���+��#�����"�7��\�L��%�� ��J=d��	�޽�@����Dp��14��B�>����_"�DMnWҋ�*���@���k��N&#�ʈ[�ѿxp>]��f2�)���DY}e�3��2)zQ��x"Ϟ����&@>խ^*�]L�TPX�ſ���~�w��łR�Wo���'�v�%�=�)b�׬ H���8����Q��j�"�;
�a]���nP\bb�EL��:WȲ\6Xy�f�T�"c���{�/
���������g�=b-YZ��ؓUX.��>��T��U:!��x�f9���DHL��6��)����Ʈ�:"����F.%jp�IG�d��R�&����a\z%�~e�u-�!����)�7�Xa�JGW$����e�P��&�FGǎ^��,+�R*$��Fo� �~�	f��J���<~�M�vd{E�իW�7���Ĝ�솬w���D\�1$T�	�L?~��)J�F{�1~��O�Z+T��j&�@yR��ro�G��臥�J�d
�j�ڗ��L�NTք���0 |�Z��H>���=P�"-����\*�U�k����;����N*6�P]d��ؙ�c�Qd�`�9;� �[�Q�֐u��S��O;%N�5�B�+[��Qʤ�� ��}\�yU�����s����Z�ms���cx���"g��3
O��t8'����@x���
y5��v��g2��Z��s�A�+z=��`�6�Jۮ(������I~��%H����>�/u(��Ih��ܴ)���>E���r��7�f�7�M4��3D4%�����5���)錬�L��?*���u-��q�"/�oF�v�<ο���\���Ԩ{8�E�����)&��*K;�����@�l�)���_�6��܌p?���.�H��0�}o_�'�������Pɋ�����j}$,ژ��_����n���G.Zݽ�&�s^X�ouР��855U9jy~=�F�yV�b��z��տ���zl�a����1k�[��k�ɩq\��U��߼�R�9?��df%�����5��uf�իWB�➞�x���#<k8���8e%%=�0����p4Z�:�B{�5?l���$'�[�&j��;��!i?��^���H$M��p	����A*T�â҈Q�mT�z|��GpW��L%����N�y'��͚'Tu���oJo��)�=:�C���Lׇ���M���,>4����~!����٨r@�@����|��}��?3=r�����/�����dYe�|�ʓ��C�O��	��������Ǡ����6�vj��㗷�5�{��Ւ؋�I-#L2A�ɡyMPr�gFщ��Pr���ʶ�ӂ�d��������?�N�!W��""��x�O �^&���|�v�J<�u�l�r��F9C��#����g|�M�۵�#�:��M����/���|d�����LÌ�|o�krW�w���z��>�:\����Nx;�TV�8�@<~�,�y|o?v�GF��������U����'�ċ]�Q���>3� 3���7�@�o��̟���D��Eb��ŕ7g��>D���@@P��X����E��`�V����ʛ6������63����C�7�cf@C�jt2՝#p��X ��x7ٳ~c7��1��W?��r16ˆ���3o�?�m�ZKL��*�����U��{ITm1b+����k���]|���Sp�� ��~�9�ؾ\�׌g0�������;�%����	g�UE��f�X��7��}�k`8��z%��ǧ�����r�rm���ݹ�oy��/�V+8�G�F}-7�0��~�;� ߯�V|a��4�+�z����X��M�'�c d|��[8�M�/��2�� Zெ���RN���Cq�!�/�<=Q4���.d�qOqv��+�>�_���>��R>�D~�$���1�GE,h��MP�����O��wl1���Z�3�i�� � f������V����y�?z�Z�U��\h��т�r�f7e�������u���q�[�5���O	W^^��a-�X�V�A*?�^q$.&F�3n�Vl-����d���#Q6�N��1�he�g�7�ǅQO�q���NЀ8��Y�;���69�n��z�ZQ>���!́G:^/���5�J�~nz��H|f3�mw޴��dSP|zc���KZ��m/����V����C��Z��A�b@@3	e���7"NɎ�J�˅��5�:�f_��߹Ɲ��5�w|��Jf�bW'Y�9ب�'�εz'����PΏ�z�d��74YM�*�:�܋�GG��"��+��mx2{��P�\̤�&H�4�"KS=�Ye�;�CIE6��ƴ���ҵ(D��C��H��JM+�e��:��+xݦX��9OL����"-f��@gBO?P�$����o0��"���������u���-)��wPi�ym�OТ���E%�Oa�p`A8>��	A�	~��7��P(�N�W�A�z�71�=��`6X�w2�f�BO��*	���Ϩֻ���]y#%.� ���VH�g��>,�|,V�uU� �[���P�_�eL�_��Cv^�h>�&z+��C#o)&�\[:o�3�6յ[XR����7:�5�=�ES��'�?[��`�Y���ܻ/����������g6 �52zL���^[��i�SW _�ݞ�O<���32?�8�p�&��D�&�щ�|j�scrv{@������QL���y�@Cu��G����ϿJ�/���o�)o�Y����>r����d���9�1�>�v��� j�����'�1�I��B3��Z;�?��@���m\�>����~J���%S1$���H3O���Z���#r�j��5*
��� w����V�.@�m����HVO����s�'�x��y{���=^r��Gj�U�G�"��}��Vv_I
�B��T�iv�����V�kQ��l�?E��i�[��QM0"�����1��̬�{3ѧ�\OaI�dl�$J�0��k���'B�a�' 4��))�)���]�X�)��w�߲��ON�|�@��?��Ly8C$IM�T�c1x|�3 �K5Q/[��N�����{��<v�%�uq�]]�o�܀���++�q�~$\~#!)����cO���홠�m)ҧҝWؿf�"B��6k��P��րχ�1��Wi͟�o]����-� ^ׂ=HT�2���^Ȗ�U������˼��ݰ�-.|l�=/�(59z�oJ���pY�ބ��������o]�(ص'3��ֺ����}�IB�RJ�Ѣ���52`zhH�TL�H��~�A�d��4�+t��+ی	XմT���B���[��\���cn�+u��mqwW��R���.��M�zg��4� �E��'�����l��Mtm~P�G�+����v���L��=�a}[����	SN���c�/��#�ӊ�y9����[-^�'�B�c�rNVc����xM[��%��!���.�7��3S���ӥtr	�����&#��=>VK\%���T����ƞ�w���W핖�E���P`�zHUȗ��!qK�C�(f7�Х߮+���9�a{?�B.��Т�@ѐ����U�2����uv*n�T���gJ��)��,�Σ�3,׸�2��;�ds�V�_>����`J�������w�7�j�e���>,�z�����+���N��4�(�z��I]f�S ������r�ʽ	쉶�i��]�i�댲�����rϙo�=�m�e�&#h���|�|�$�B}u&K�� ��٧B�뽖��'9u���ڕ#��s��r���]ɓ�����>"j�NQQS���Ŗ'K�V澷���tI�kv|�(>C������%$'��Sꞡ����J󐇛�z�N�	Ʊ�<K�ڼs����3N�'v������ַ����^�Y i�����H�`�����G�b�k:�:��}����\�"@�]�z�iM1�mH4��3�!��,k�Ԉ����b�_ִ��+�<7?�XCtޤ�ω0�5.��l"x�F��C�C���Lm�X̢���2w�8���i��^��>֬a6z-b�R8��d�gZ��Z��z���Q�jH��5���v8镳2ښj��֋RR�M����ץ��J�yp¶�{֮�^�b �.���7 ���O=�t����D��F��5b0G�$���y|�ܠ.-��U}����Y�[¨G��Y�bHz��K��f?M5�Y\��K��f'�������j�q p��C��H��v��K��j�6�Q��C�f��qP��Sm�d,�.�:ʘXs�F ���;�ؒ��ҽt��L�����)�M���6[��h�ëۿ���,\��c_��l.<�?�N�<��̃Tb�1�ǒ����ɂ�q1/���J䱇��tͻ�{�>c��Xr�X$˝ӌo7/on	�7[�� ߫����x��8�@��ZѷOƸ'�l7��`vR��G�P�5@f@��2�D�'6��X0�m�"O���R=Ǿe��R>:i�5�|\�r�%C���LY���y����m�-S[�V^e�*s-���_�j�f�Dآ8{B�˶���T��ĪϷZZO��k����]��M��*��� �wl��nc����5�JO������$����6�(�M+z�҂V�";���Ϡ��W�p/�d�?/�R
��ʿ��^�pH��+��*���5zd6K�	��iRe8�$l�Y�pD�O��"p#�|��CA����#T��1�C�)V��(1��Z7�upߙe��Ρ
Ł��1�o�shP����p�Gkmkjzm�z�����6��V�������5��:�3��j0���G!�1�����Ă����>�����V��������BN���K�C9�F�CS��j'�YD�����=U��z�*�o��f���.�[B�9L�~�#7�#���:�ܽu��Sr)���go���w���h�v�V�)xsʿfr�P���u�#O��v��5(��G�4~[ЪK�҄�T��xu�E�wWM��|6�R fs��)"�E�c�֏���_�Y[/�4&�|)ryef�޴��L�=d�`��A��=X�b�M6�W'>�n�>j64���P��@}�L��&��!�%t���
�}�����_C�Nq��q]G�T�G���{f��l	�b"��jc�Z籟�R'6��&|���>)*�zJ=��p/Ȩ�7���fKve���L�"�r������<.�Z{��ؑ�IR���A���>l��������6�% �r'����6�F�Lw�gm��<8=SQT�ez��\���QY���u/�Y�>;^��\Y��<�Vd^������4��*@�<u�4�[��	��U�1Z�pĺ��b�N)2uXF�]3e��Hm��=(��V/�f�n-ߔ��������n��6��:�r:����]ss�ޯ�o\m�'"OM{{�U��#����~!���t��%#�>�&�涘 �"��%�ٞ�������IZW�o@�_���XԹ�x� �1	�׹�ܼ��!���N; �*��A�>�j�B�<�9zۦ����+ut�>ɘ
۽o�-��q�����*�Dŷ�b��@+��)��K��y�[�/GQ׈WRS���x#�Ej��Z��㏻�����r��]Ex"#�"*�S�N�-�Ddk��g�#j�Ï��P���s���\�-���˴'ּ��tЇk/0���6�U��eA��>�s���?�9*�ϡ���;rh�.jz�{n���,�#�|��l�c5	A�o�
������67���e������7�p�	Uz�2;��I���,Y�=\WO�YEc�ײ�ȥ�C'4��X(��f��k�dT�E)��:r�i�nX�V��^�s�Q�����Hl=q�wz=Qk�t�
�z�P>�EA���:+�U��a�о�}��ﰠ���-�@$�����\��<9��%�$�s
��+���P��,�R�ʝ2\��0�}�J�f��Ipꨣ7��x�@�؉Y�������g�o߰��ի�S��hV��Y��=bZ�{�i�t�&F�K�/�u���t�3&��\b����V���W�fN8z�$C������#~͓�\��

O�~���<E/]	DY��P�<���d8i�H�|E���m��-A6唦Ӻz�^w��y0.��@�~��5h�`�@���VՍ��/�/6R博�����y׋x��#�3 ��͌���Vz�����#�}���4;�!c�R�TD)�.����	��-aL�g�^= "�y[��I	�Ҝy(+�z����d�Cl{Ֆ�F(�/_�7;r4M���$$��3h���1��L<u˧(t�oe@��a���ٝ��MZ�F��A�
ݗ�{�R�W�X}Ƙg�j��R�u��k�1M�A�ޯ�0_?Øz!1c�V�"���v)��?z0������oЀ?l00���'R�mҔ5H[���*`�~��>lv4G�1q�7L�叙(v����3_�o���u|��?~t,ț}C_, �sG핻��g\,ʎ��s�ؗ�8��p�r��&o��2/�u��'���o�q�T:zY��f�_��c���kN�V(��ijT�5��'�"4 Q��*���\�l�B�y6�^��#EV�H¯j�����g�Y՞���U��;����\��<�����]'q����yĩ����݌gsq�(�`�J���qM�MI,�h�N�ؗnD�Y�ln^��(�i�����PBXX݃\���b9����I��ӫ|$׶K&�3�\ba����#e*��7Vk*-5m2 +��}����fc>����U*f`6Y�"����)��6�Z
툅ו��/T0�0��>G:	z7h08%�Զ�)?�r���{�S	j��LM� 4?HW���`_h�s��I@��Qs���i1sk�Y�Y&\��}���2 ��(�pRDl�܋�d��r@6E�)���7!d����r�S#x<N��.ܽJ����0٨���j�-8]mt�(�Th�Nbn������~���}vP��-����%�Y�%]�� ��tg#�ܥ�-���Q	.բi��>߫���Z�h�d� vW�y"nrʱ��g��x�ku���X��a��%��Ӄ���%�ЁXTV ƇP�U�Z���3��h��얃�����f5��	_�E�V�t2�P{�^�v)��X�?ȷ=�r
뫷[,@ Y�; �T���޴Gդ%��Ѐ�;qУ Z�+ܓ}4J6vP.;9LAS#.S%��[����ljA�j�y��q]D�)�k]U�������79����|`���J:��}n�r��.ט��[L��CĆc�Fu�;�+f���"��aX�^�� �+��̩ʻ�'�� �g�8�4f�y˶�t�?�c�|�.i��(r�
��d6Y�܂�]��S)!���[d��M����p�ʖN=K7�Y
�8W+�n��%yLz��:�ϝ�����I�(��Z�$= ��k����m�q����X�1��r��ͨ����,���q�?��ȓǜ	Ks�|� Y����8��\Ir���U��J�3$�YЬ��$����('^����o�(�K�I]����x9��-��-&�e�J��[�������J�))���Z�0�+P�}��.��f@-���Gg��"�^HdVk��Y�|X�f��$k� �i;�Mk��OGj �9��ǋ Ӌ�%|i�\�UW$�?Yt����aZ�>�4p̕x�f�asҜ+��|t|)M�[B�q���o�|�Sļ��T/2�j�\}*���`RO/J�f%1���͛@��;�8����*����Ý=��wg�u�s1����f��Aɢ�n���.�IO����@����e�i3�e�ZX�����,,����%�cҦ�<��Hhn�In�d9�6`�z#�؂%�'È�-�F�7��ʫ/:��@��q�)�8/Ib�-(��:�J��_�o����K�#�!�uJ/��A`��vvIj��S���%�+Uc~Evj��d��c��ꌵ��>�t��2�����`����<Q0����`j�{|l�����zba]�E��!�:=�νSdKy�o�/:,�Ald 9�돦ٸnG��;k�� ��l���P���t��$����y!r�KƐb�yi�5���ю"��	a0�p8�u�ԡ���p���T�0��#�'��
��<K1=9��/<MJ��/\��^ �����OYn��o�����"v���[����Y���ef�\�u�}�l�A12�i�.-�t�g#B,ފ�pOdn%�ؓ�"u?������k��a�1���B�*�+���ð���
au�Y��|��w�5Tu��T]f�}�Jº�- ��N��L���/Tz�њk�^���O�{�%e���p�S)BH;% �<ۭ`5�B�S ����Q������mx�^ǉ�����E�3���F5�*�C}r����bC"�Zs'lȁq�LC/['��?+�u�0���Xn�:?�u���զ�Y�S\N'���e�2�Yv���F��n><^}���O3�Z��]��	���+'}�G�5��{p3>�Z�&{g�Z���|���mJ��^/�p;5!�
%�}�g�`�"�7��HgkÃ�D��Zk=��Zh}��OO�˫NL|T�뿙���������8y��+��.����k����u��AK�ˮw���B�3�t�y&�����8n����ϛ�U�&�����ǢN:��%xN	�n�%Í �1VӬ\�� Q_9������U�O�m_NGӏ�[�vB��mJ�^��@Ң�K�X�1����!��O�B�S���"P4��Z�O�Vf��R��{���*����ߢф�
�==���F��&j��;7X���#3�S���UK����gS��%yf��$CѦ�7����������\ � �W����ޙ�������A���c��T��z���_�vK��]ݐ���:��n����Y�(���k����sJ�rͲ�����t��j*MJ\\��[����׸�^�.|��
��6xic�����p�#kp����][�V�H|�^��]qau��R�-��nUWO�P5o�#o�zm�.P���Y�Թgz�Ɏ�j�_a�Z1��׽����u@v�@��������H��ck��W.~;K+Y�/�l��3]jg�=�S$2�D�:��+�I'[����H��S1@�ѱ�k#�y���7A� �@kbN�6��:���ϫI�F(��{K�q�ڵ��)vI�6>�<�%�?�'=�cz��܌�p 1�<c����l�K����L�Abꑁc�'[w
��5q�D�)�E(U��像�[3p��|b&�~'�r�GQ�g�{O_4��ċ��f��P䰿IS��W��ȱ{M�Cʟ~D3K�0�)ּ{ȍ��,:�'���g�Y�rzR��ԇ�6┍8�A���z���:����mJ�&����Zʺ�B~۪���=L:<*I�z "0�"g���oO�~-ɥfw�csQ3�DhOʰ>��KGX�`��P���ZY��m>re�lÏgD4�7,����0oee�Z޹Mw�2�q�,N#4���6�3+�����O;���1(���)��~v�C�UL�Cj��gN>�ݾ��}w��)y^���QD��L��s����D�z��	�������rS|m�flC��_9�B]�+��Y���&���+r��&8��ϫ�}q�q��Ag��a��3�⛱Z(S�����r��p�9e�|M`�@;`�?����B�Dg�w.�A2�d�,'�J	�e�D*��wbT*45��z�`�C�{ WSRЉ1k�b�#��zN֨j�g�R�ȮR� X��=5�ed�;� �n�?:����=x+�AU�h���ˤ?���a6��7�*���!o�lv0�ۧ
0�)V{�xn����%���?�.xbtӛ� 
%.}sAN��k�!������p^^���Į��EYC���j���R�7Z<?��:���QK#3��-c���}Ѐ�rM%6ȑk�� 7M�����0HR�`(�[�"�#���-�Ε%5������YU�K<��n���,ֳ�|zp�\X�����6��jOj��R_�/$X� ����eA�D'//<���$��l�#��ݳ����C��A�C#D�������?�qD[�A�����xK��k��1�O�է�̲��Ջ�}އQ�e.Q:�HJ�Lx�|`������oT%{��C˴>����%���6�Ꞇ<eY/μK@����o�&ce������X��i�,	m��k��}^�h1s�K�n�>��М�I�]k>_�$���y��&Zp�;��#�v�o�+�����p��0�`�=B����������qH]RK]��_>O@]��Y�֦M�ȱEN�r<qi�:��Z i Q6��lX�%`;np(j�3�M�����/ii% ����il�Z��b9��8�f=�4hD�����<���:����Ma���!a��W��(�л��gV&NEs�ΏZg���Ż�|�˃�шj<�:�U��1I�aH�퟿,���Ԏ���"��N��w�?���\�h�y`��Lf#��m�*�Q�^��ngq8K4/��������t���;���
��X>Q��h��JZ@&�y@ܯ������ӆ@�H\\���%'6���5'������)�D$1����!�v����=�IH�D�h���҃����B��q�B;rQR�H��=c��EƤDdo�Hz�.Q����\�A��N�[{�¯i�۞�;��(���E��f}��vL�^� �0$���!�z$ �O!�Օʫ�T�,
�Y
C^��wۀ���O� ^�e�e��b��/���m���l�l��μQ�L�e��Ņ�ZS�ev��Zq=���nR���x���ݭ}�,����� '�R���CUPb�ã�X��5�ئ7���]�ρ��m#=0s���`�������������s) �o�K 2��}P���� &i:�����j�p��(�媆m��m�^���̃�O�b(OB!�3�qV�] ��.*�� :����G|n	����h�I{ɻkn(��5�mr��i�v�����W`��,��cR�>*�k�'G�ڀ{��w1�r�kʟB3�s=��*w����� d���������
�t�y;mh����d]��ٸ��������-Q�M�Q1WH	�A�x����;�#E,�eDD��5��z��rVX�������B��ܛ'�'����w��V���}*�:io#֕���Z�A&���c�LV������}������.;�/С��K�}�Tr�8�.��7��M�L��(����'�vC|��#}T%�J��9a��H�%��{忥Z�Ԉ�Ă���c��ּ�[����	�`�Õ��rb`�^�4m5���&:�^���������7?�76�%G�[�m���i\h����X/0�E�Ը��D���y̩�ܻ�J�3:�2#�> ��Y���Z���j;DW����7�q��-��N�'c]x 8
��a:X !�(K�{̀,U�K9|ZI�$��O���8)��"��0�o��po~���c>$���E�H�����-p��^w���~{A�#N����ö���󢉭&&q/�����<�Q��u����C6���*HM�:��T��]Zx�<�h>���1F��`)��T�ڋ�Y�o�^|�u�I��<��ܰ�D^d�@>����c!�ί����r���Y:��cʒ��{�˔�=D��X�������T�[}�R=�" ^���bV�Y��~Xm����RD�0G��O���ަ�9�� �i��ვ�@׉S�n<���N������҄���/�U�ИD�NiȌ�}d�Ɋ_|,��1UL��@tF;'.��_��涴��8(Vz֭׊8u�<ꨅ�댙�Xq<n��Z�[0�XX؜�c��<8��V�c���w�*�R�@���2���~" _�
l8 ���_�%h�c �Hu��K����LL��
x��L��9�>?G]�xϒ��^X�X�B��W[<yF��	��*���I�����pߡW��Q��i�@���#�h��3��~�8�����P�jP���1ſg���Ʀ�򫝾%V�G���$�-��sӬOM7�p�q�����jL��>��AY
��?��z��"H����(on��#�|'���c	3��bL|�4ڬ>?�5S�eQ4��UTT�A��~��l��w]�z��'��mʈ]#��!~p�L�a�,��+�س��kޒ����V&�ꟀGiL�*�{拈�a�?���F�l�c�2��敟J����[��>:<�iR�&�P��e����4���99����&�0��}����������t�º�����T�Uʆ�MK�${u�Ø��@`�1�{J��U�&Z��٧�-�V�.ϳ��~���A����LNJ���M�M�X�1W�V�x�����k�Ap�có"u~��u��@7�M�,������j� }������s���=�Ԣ�28�#f� ��������J�9x�@�ğ��P�[���\�3i��hqr�2��wx���l~l�*KV�{���c/��,��F_�4�\�ތ.0�,��U����8%��I6�^��U��>�|�G��r����S�l�N�x���Fh��|�1p�*��X^�s�Q񊕈�=����	����\b!c[�����{���XU��2��v[�65�Y,����z|M�у��������`��p]���p�=�\!v�7��<"�C��}�<��ܐ�v�X�:���s��;���4�33�z�Չ�_�B�����=8<�1�}����6@���Y��x� �D-K��3����ދ���˵��Q����"`������ƣ�!��LK�C���{"O�m�҇���j��	x]�~wI�F���O�|�wן]�|!����+v����$ro��5��/���]
yCr{`���Y�I��9�˳��W^����0���|��2�o9�	�����D�B���T���7��iK_�t#�Kt��1{n�-E�O�Au9h���,W7/y��'�/=�����;�֋fB��u�,Ά�v�8��0Jy�T��ޅx|������'�q���r�IM����������*��t����}C	��I�H��[�~?���3њ��Q�Y�'�<��� �v�:go��W+��V�¸�<[JyZϥ���_Y�H�m�|fq9�b�0]�9Cȗ@�rUk��wi��U��SPý�����'�蛥=�;�B�		��x(��}	)�W���u��]�F��Y�k4���V|fu�}|5�ה�y3�sk�B������ ����0>���Ծ�v"a�󷫼��.-����f�]�u�C�����?�tS�
_����[�Y/G&�Yq����cPa�TA2�Ǫ�����ڕ��?�|���jT���.p�0弛5�P���q�9�[o�N̟��(Έ����~����=��3^���ꭙ�.�АKb"�T���a��w�����Ņ%;�\�LYB��"L�i��L潧Z�o�2o��8��|�*�ǁ�����n{d��&����}VV"����*�"j���+�����>�$XZV��s�?�96>��ߗ�2Um��]�:�,�%����������z�����c�/"*����+�:��(�� ���w柽�����y�tu��%��������v�����
�X���tp�[�'����7������n��:�PO���}+������x����Ľ�2��>�ۖ�ou!c�v�����{�!|�������M6�q�������Tj�Ԥg�Gm�������j�އ������CBZB��������K����n�z������l�>g�Z�z�}�g7Hg.��ұi�ӐHd���م}���=c�ՋE~�),ȫ]�-�W�u�NN��u��"8�h
��y}@���G�������X����IXO��JSF \�8�o��Jr,���O����0��U(�@��y��^s�T.�s�n��/S1�Svھ,gsqÛ�y{6��� ;�r���������c������X3�9��s��'�p�1p����36:��9:�F~n�jd���*�qWo&��nWp��]��S�+3��L��	�=|��]�>�-��M��]o�~Y�U�\2��)G����"��`���d��=�`oc����+Wc��O`|�<o��U'�!�� ��c}a��\�(��,3�g+h=���ɨ�L�I�w���(�k2�A��(b�FEj"�&T݌����c���F�ᱣ�cC��+K��4#�� b0nK#65���Ǝ����z���Ȟ�0����o^5獽C#,�¶�bP?	�j�R6����Ց�s�ҟ��4ᒐ�D��CJ*Xo�k����%�<$��Ƹ��+��(O�s�j6$�U�F>��.A�\s{�7%��yy�(�)l�=�B�=���=���y{�e-AxrG0�Q�����k�*��a^�]��f{��砗�ܪ~H_j�l����lg%7��oʠN�����]��~�zywhs�*F7�:��wh�����d� �ϥp���Dk�5w�I���N��N��N`�\�n/�,�-V�P��6�42���&���o;�	�GY��t;�y8#K�8�	�a���.��&ێ�_��<�ir�׊]��;��\!3��z�l���ptG��)rI��֢A
�
~g��VBn�B�F:�L?�/93�$;�����dN���@ܿ'G�5��7c�=Mln��g�Gw��Ǽ�����M^����S���ɴ$�+i<.x�C��u{��:p6� BC]��LBFBY���pa����y{ȅԿM�]5����[Ն�M�������4�#g���X�U�fg-ߞjܞ�8[/�A��D�樉�$l�̐ۈ�m���r�~�����������6�nd�/u�z��߫Ȍ��6?�
A�['4��D'���e\�l�:`��܂�����Dl����|~p������D��[�l퀻rff]�ן
l-���s�`*�����uM���2��I'��$R	C`��d������֣7�_*`@�6GQ�e�!i4'_6��(d�֓96��;H���S��N.] $�	2'�@��4�18O�W�n��T�	0}XNB0_��@��]0�Id�n�`-�o0�`Q���+��J��U<<<��)H�Ŕ�uY[��fw�}��������R�Ep�D��).��}���,+)=D ��v>�b
m,�p�'kp&h�-�4�0G����S�hmW����>��]U�wb�eb�����K�Vפ���{��Z��ͼC^�H��"i�}�$�;t[Zc�u���<˨���ͣ�Tkzkw���'�{!D�-�ďS�ꪂ9��D{t����o�9�̊IΤ���[Xj��Nv�d����x�۷�]�ɷ�	L��K��GX߶�¢��r�M
��[@tM�,"�-��a۵?�!�R��Hd�yو�:WO��8[��0�/S���ъ�,�dE��T�*���YBrYllB�h�./o���Kt���ۣ�-���T9x���'~��i��:e�K,� `�0��0�tȞ7=��m�vo~����O��,쁙QUkc&�S��E��������=YHR�
���g�n�lgoP�w�[�@�ɲ�B�������Ê�%�(��6��=�k��jg�V�l��K����JY�H�{�pp���C���2�"m��a�?w>i�xq��D� �u�'UB���ձ�L)�|�W�Qgs+��+Ԛ�L7M�ə�yD��,��/-�fy��O�|��d5#[3h�D:��U������	��+m�@,(�ѫ�?q�O��y���E�30/ �������BWS�Kq�#�07fhfUQ[Aǟ빧��7Z=��Y~U����IԷgaA�x��w�9=���-��w���FD ·2��4��so����)B5�R����	�'�cӉk����3�<p-��|k�=_x#�Վ��7��Tٳ����j����o�ShT���@_$B���|�06&����Y���#���>	�t���0���n��>���O�6�Wa�0�-T<
�(��}gg�ӵ�C������H�%|��j�ɿW�P{���N��o�ה�<�;��u�}_�j�]]���{�:��l��ν���F�׮�ec>���mӢ�O"gy5K>�}�`�|L��	��0�s^q����^^K��LY����Zyj�]|�O�^�w��v1q��'k���y�Qo�v�s�n+K��МI� �DQugd�F�����"��oBh�9�M���UR;�j2.kԷ8E�;p#ր]�.T�j0��E ���}Y��'[�Q��P���A?�G%P���c!�{`�nwP��1�&���{t׈����)��E�/O^֏`�?&�>7M�ea�y���J?6\��[�e�2�,�H ��5�;]�����/_6�,��ڮ)J}���*'6��س���N>�����0%Lz4ʙW�O�ȵ�>��v��d�@?B"����4�|�uӏk���6�b�hw�$[@�y�}�g7M}v�,V�����tQNd��?�!�ct5�w'��ZX4�4On�45��ka���@�Z�#γü�á�~���Ey4҅a,Zn�xQ�6.WA��?��L�
�d�A$Ғhv�� �uO�3y��9���L����_��Ĳ��F����=��ҧg&-�03����K�ӎ��| +Jq)ۨ��
X�u����Ϟu�hV]���ă������1\�Wl��@�!v�)m���B�J) "vMu#Xq?����l�fFZT�;����)B�"�����)}$i!�!Ao �����7�l�R;�k6[ݠy�Y�8��VEV^z��i�����7�U�@L�ټ�� W��.p�:���p���J��K����]|�P
~��N;(x `�1�ۊ������6b�;;��S�Mr���N�p}b�%N	�M��	��	�&��b���78��n0��=�;i��"u.�����e� '�[lR�D�R�a�F�zr��9p�����ד��U?K����>��v�:,���B���{b@��m��,�?Z�\Sߑ52C���� �ʼAc�8�F8i{|�X�$�U��d�*Rx�\�cY�z˅�ADozcǼ~;{"j��Ʌ\�8s�����7�K_3�m�q�b ��syXOl��
��!t����`�����#ܚ�/:�~s�^�����6�������wM}�W���+�L�_ฟ�DK��I�ڝ�2�ǃ�nb�2��P�����嘆'�_8�~���*�G͆�FYȸr��Z���p׳ċ����٭��C�8�?�2D>ڷ��]i��V7�������U`*�Ɖ�b=�->X<c�ւ�ر����p%���ʷ�kPW��\���1v$)���wj���G�����yu��ـ\BЕS�(UM����b�Xzz�7Ooiؽ��!$_�n��@.�"�X�\x8|P�:^$H�Z�����w��� �;���
���\���R%CZ�`X��-�~��{eu1�F}�H/1��z&%G���uh�����b,ZF%�`�Ob<E�/�e=�J�����������Nͫ�;߂��ƞ��+�߃sUԽ��K��1e�v�����"A��D��L	���(�j*P�T���m��d��P�}r�YFY�#D��~\��)I�tFU��slF#�`��m�h�Hx�^�(ke_�"��g��o�WVĽ^.��0�"9��7� �-�H�Y���$�*â���{.(�M6��gv��2t_�3?'����DG@��ڸ�j���Ȕ�m���S�y�Y�O�շ1�D�ٸ�A\m�>�K=�� �/s�r�����/��j$ow��:���0��-
�,6�&I�+ �-ߦ��уԮ�? m
~�F'��� ��i�Di���Ĭk~�{�7��O��/� _��-��;��z)�fu�	����H;�9,��	�{����Y��.�����! +&�f#ؕ�����9�Z~�����2Hfd��_��L瞂�
k߀��(-�5��B����]ٗ^������$��n.���W����H�<�������?3/k?`	h�L�����Pey]�UN���N� ��vGO�c�p{��@^\gȻ���&�oU9ʮH>NIj���`"����j��΄��	kňj��ͲǼ�S��$� ��q���*T��oŶ�ZT�@e����S�蔄�cPh����vnET���J����9���VX�M��[�J/:�ՠ�J�w���!=���#*Z����ץ�.];Olf�7�!�l-�pC� Ġ\��C$���m��g�c���c�7K'ֺ��R=F)�PN����:}���O�,a�TvW�UN~�%�F�����{�p��:�My$�FI)f��p��w�-$!����ɧ}��̊�à���(���E�AF���N�ICc�3|��"-;4fC�G�a���s$�㺳�s3�|ͯxݶ�u[�A��܏���sւ��z�'��c�Ľ�]�d"�m�.�IRS��]����C���������^�.Wն�2)7�yp�L_c��A��_��ԇ���G��PB�?��پ�#��s�9�^���[͇U�6~�m�R'B	hJ|~0I��
{� 5�k�h���"��C�#拧'
>i~L�
��z�>ilM�?��+���I���h?�!���7S����R�6�'nK>4�IF/I�gݹfl%`:�f�T<�W��.�q�::r��"ϛ����PU~���P�W����9��3Ő���f7\U}��h&�x�S����N����v
�y��;�g^۠�,yl��`���ʸv�dK�s;�h���������K�Z�#_�=���I��|Ƅ�N�1�|uC�L�5��ҀH�@5"F�H��DZ�{���9��h��,V,�}]E�y:E��������7�y�'�WB������OZ2���˲3R��B�/o��W��|jǝ6�1��<Y5��.����m���P5Xt�����p/�{�d��TWs~[c3�I�"�lUM�����Y�B�99� �'�[������V:�q�`�\���08�A��Lr1 ���R��{���ueTٮd��a��w�Q�{�<�a�0�zq6�R���ն�=��֊��PM+,��&QE)A��L���][l7g^�4�O�qC�ダ���*�ߥ�������n�V��A���Ő��ެ/�5D|a�_����L��8�m��$�x�d;�yh�]W�t��r�<A;��ߺ�ʧ"M����p��&W�݊����_
 ���G����a2�f(��-�2�z��t�f�.�_���r�4p��u4�/$Fo`z�S�U@��B���U�&ig�y4 P�n�_�u�Qc�W=n/9�h;�6��Ah��X1Ga��M��]�����^�)��kWH�Rl23YI�]��_�)�q�A�-�3��n4W�	O����z'}ї���FV@�]�F��1�Ms+ �<�����y���E.�&s�{�b4���p����x�����n��ǰ��A���5��oY�@�O�/-[vP�tҧZEt~�-F�3�Yz���@����_݊֩���Nt8rK���s-92)j��.�������%���<4����j)7B�k�\w�o�y)EQ�S��o/b�4����fYT��k��E:�IY58\�����|Jn����`M�G�������2�(Mb�ț�G|���F0�ϳX)u��_���
��;�;:�oN��|N�R�6K����w�ܤ���=V ��s"#S���hm?�~�B�c���s-�M
�0X�A	Y�F�#�6�I�T^s~��N���$�}� ��e�Q�%
�߈���}
���0&]l��_��o�ѯ��1�* �1b�X��u%ō���90���?Rwf#)��S%ʔFbڡ'�Fm~�==fb�0��PMᯡ�'㷹��H��F�IE�탓|�fw�[�>X�[ۼK&��`�
Y������۵y���
SMq��v��eo]��=qPw�{��Ğ<>.��/
Rf�v��vms�����*�%ƥF|el0\_�X+��-��Z����:꥝�˸�E���f˾@�7�%ˬ������h
F�U�D��\��^����l�`Q�l���%u���lAۦ��F����}�>��~�;KL8������ oto�*}��-���@��A�vm��m���}玏���w���n�K��)	x/Pëg�u�q������hB�����b��w��*y�\�ٟ��)(3!չfSƄ�u:�j"�� h�?��W(x�|uz���w����C'�)B�``oݺWc��X���߳��<���������P�
���=��/_~���F�]�[�CiV[j/��u\�{��3X�bd��.cP�R3bM��V��K�6�l&�>W.�a���wj�1�ֲ�����LP���f�vt��{(���aHr(_��Z,�9'E؝j̀��і~k��t�+�89��*Z֙~� ��͌@��Xo0��E��X_�������D'ڼ9��c�
C���ˮ��M�ޫr� �C'y�M�1����i������f�	�����7&0��{p3�L�)5a�wu�g����3H	�!��?gҘ(�q`�R�ɇ�5�27|���)Z��P�bp�&4'�V����C�x�/�5��lX��gS�`W���Lz��
6��bQ �4�z�T�����@,��TLg����[�z�PD��%D�%f����ڵ瘀n0\+g��<c�l�������%�7�~N��A(351d���.���)Ӂl��DaA�/����Oy�2��1ƾ,i��2*�s�W.KW;%3x���0ơҽ���A�%�O���TdG6Xs��X�H�,,���ڂh���v+�!��l��e&�%X��~�_��� ������>�5���om����n�%4Ja�P���R##d�6�jG�"*�$��q��?�~F�a�=��wB��X����GK�(������j{��e+�:��xV$��i��R_���w�]2 ;�d����;d���\���[�]�u#.�m����>��ʇ�I�PQ���5{�[T���=i^�KٕP��W*@c�:���mU]6�}�ۮc�i!�W!��lB��C�3=������ǒ��O%�����m�vL�ؑlWG����7S��^����3����)|�Yh9�c��$���[�&P-�u;ݺ�7�R.��E9�@N�� ��L̃3ϧKU�:�����3���N�a5�'�"(�e����OL�����H:>Ó~��[[��f�Uٷ��7��H�Ѐ�G�<���▙�Q6u����p��2�'u8��1�;�����f��e;��p٧$7�hv(ӈ�X��^1��?��:-,��"*U���Y�u�ܐ���fm�Et���}@�T�U	��|*~Y�A$,s����lGf��t�j�u�~��\I���Kt��-En�:�'��\�����c����m��J��ã���wM�u>�]�2(J���䜷��4)�u?���EZW3�]���W������_t���eQT����������}���c��ټ�uؾ×w?��#��j��;<\��({����l|]�����/��a�*w�^�ႇW`�H{�1�4_��0 b	�?V���I��#O�u���}��F7��^ui�����
8�T������hIy��Ke�mQt�_/P1���Q�;���j���K����}�n��X cCㄮ;�(��)D��cSr���%r�)�	S��S*Q�mMd<�����׹q8���q�r�6xx�]��z�A�����7���8
Z�������[k(��_��W�k~b�f��+�,>�2�hWU��_h������E'u���Ht��u�2����7n����y�Hf����Hbݶ_#�F0�o~�}��i'���~`Ct@[�Y<R}���o��u�����2��	o��䩔���+�qjޮ���X��๶9CjLk�3v$��L�s���fWYy��<M�oT��n�I�6V���m�nş�	qMvS(��g{.P�/��Q���?��#�%zN�K�����!y=K��q>��1�<���}:}QR��X����ѷ�����I`b�_�"h�"MW�JX�8#fd&�o[�M'L�bR>��EQr��w�B�,��r3ʁ��ugv��^�)��:�b|ڗ�Z��'�@�1t#;aF���ê`^��P�D�����8�l�2�]HqWa�ňQ��h*�� Wzm<��<yd�
���S9XKɕ^P � ������C�Q�����`4[0 e�o�hj�n9R������v�Q�"���8��}�auT=;wd�_@GM~��W�3���^����<�}G�%�מ��YO;V)Nj� �����AqPڥ��^�%��9�3.)3`MH�������A�r_(Ťy��-c����������K��bN��� ��� �Ή�XG����g�垉��=IJ�:�D��r�� #���1����<<�������2 B��_D�9y��+x��CG�9���X���͝ɲ�<���_���ۻ�C>sb�P�9�bp��j�'f��Q����Ic^�z�����{0��Χ8�fU��҄7ߧُ^.�~p��\=�~�3�O)t|$��FMDfV�!yn�M_��P��C�'���w�x���u�k����(ll:�@^o�z���O��6Ul���)�g��W׺d��h@\�"�@��@d�{F�\�~�h�z�`��(8����@n�~�Q���M����G�q�\�JBr���C���~*�?+�� �uW��g~p�&�sh��_Z,�`������K�W�h��C�՜�|��;��ěg܁+��jQEU��r�Y������^j�<>�2���݈��~h
I�V&� "SRE�g�%��Gm���a���Q~�0���+�!�����K� y艡�$�YG3�P�{��>tdGSC�p�;)7�;iGE������5{50�@��7��hG�_����{���!������1W��w���>�|н�&RWJd	eJM���d�?��K T9'Ņ���-�O�*x� <�-ҽ�+"��s�A.q{��r�{M�-P�	�O�y0�I�u���i�=IL�}v򢎲���	���Ɨ/�P�!�@!�?[�M㹙l#}>�`U�~�$�Lqw�G�IS��] �Spg)���A�c۴��p�@$xB�����ht1U��:@�����#�*����g��y���k�DB�+�l�kx
C�T>cqܰ�Sd��:�eB�v�i���Ƙ���O�ȟM����3��ڷ�!���J�q-&[�[��Г9��TE���i��* ���D�{T���ն#�ҕ[�@<���n�*�8��s�m�����B�2�pD�S��C�lf��a9�,�P}���C�0(E��:��ˌ���C���5��Fe����&�_z�R�e#�%�I�ք*�v�+$�S�7e��ۘgs�[lvsD�i\��6���{OO���5�\!@�Q�T-��<�7-*��n�<<���Ud�g�����)̀�V�,�P��|{>�I�f)�(��ϟK;������B��<}�1<�9���D<|�0�ؔ�'�&�1��0^(��?��.Q3��˩ӂx��=zh�2���4?&��aL��P�?�PQ��o��`�l�L���D�A �[�=D ,K�,��Ds���>@�ޣ�`R�����8Ƚ���t�=;����\�R 	�"�F���EA����<�zLY��G!#a\��
O���j�=�Ӻ~���k��~�ШΘ[a���z�OU-�jY�;${y�ѥ��1--��'_��X2)>9),�k�%�f��毷����]X�𱤫\��y�x!z��l��
��b&�y�e���L8�l�Z4f���3�D�M� �E�҉��Y(�\"ͳOz��#��ۄxԻ�����Ӵ��C���,M���<UX5�%O�ڈ�lo��UU��%
T���7��������_�y�yPZ��$����o&�WvN�%�Q/�`��O
�����U����x�S}0�so�&8 n�R؛G��mz�oOSyND�7�|�a�4ko��`�����)R�ǰIˑH3=�p����R�����ת�xmm��� -Y����� P��>`�0q��0ڒ��xo;�V���զ;�i'Pg����ÈG���[1Fw��b������%���/��!O�q�*�o���u�
��+�$�F��tH�گ 1��X������?_T�'��`eR(�ebSq�g�Z�nF�y%邾�����C&x���kU�����ܣHM���9B���i��*.�*K��s�dЖ�\q�ڍL��W�����xa�w����L�����̯��R����N��������5��s�I�X!t��fU��2@�Cm��sN�џ��X��x�*KO�3� ��Vi9N��� X��BOa!>j|c"�}&��if����5b�C6��j�ɑ���=%q1#6�˲�Ȉ�S2M5��H��8���	��?�AD���u���'�,t�&��`Y����}�:���R �W������q�<�eeG���R3�����l:���$��$ٟJ0`'�����	&�0=�ⳋ4{�@�d����&�u���.�-�/Gz��K#.�rh��",��'��Roa��?�0`+x�@�w��&��r����;D�h7�Ę�����{�I�����k��Vb����%�ט[M��7$�k7\�����A�	h ��D��F��.b�#�gu@��Gx�<PC{>uxK\�-ፎ�*�k���;އ���]+0��^��8��,�`;X�qi\��/�Q�̶
aRa�X����㍆47�Ym*��H�KW,O�zY��4�˜�H��^g���A��<��)�����J*�Vs�}:t�т὘��e���L1I�D�1y>ܤGK�V���ϩ�2�OCP��2��y��h4�1��J	qīCf��D�Fv���`�a��	pX�} �U�q!�����LZB"�$�f��?��<�8k-9���S��9GҪ�Ԝ7̠��C��p��.���6Г������=�>�p��RQ��7�g�e�:?���|"w2��h&m<3`z�q���:�B��(��c|�w�Qu~R���F�7�L�[6�C�`���<~�0f�W�#h�iy��%<2�9��L-6�u��F�pa�h����M�] ֪������i��T� �z�� ���B�coV��Z���[U�k\ub��/�HrA�ӡ){QSt��ZfP<����T��1�{�����`�/5K�<�G��"�]����,��s�c8�'�\N�pRu-�x�6�����Cc�O(�e��/ŏ8��ZD��V_ߑUD�2��E���".���$N�A�t�j�)Y �_���՝/�&�+����S	٢����g�TE`Hv's�w�c��@���K.� �M�9�Z�T	�(��g�Re������!����6
�?+'g\�d�G�par�y��T�Uz���ɚ\�T��l�Hh�h�}0�쥝��ěol��+�v}�-��rz��6={顗ƈ�+���R���!����+��}u"+�Z4�<+SV���ό��7��eI��߮hg5{ϞJ���	ZҰ�跪Ȥ�� �ݡ7����;�-��?+jɌ;�������	'\8�Y�����5%��7o�.t�~2Mp�a��mB������nd
�F����c		\|]�y�jn��&}(�6�~���O�9�H ,����5V	b/q����$��9Č'���(9�E-�;3�+n¢J4��2�q[���&�#�YˌS�/_*��Y�aø�s�����i�[rF5�[[9L����@<�y��VZ6Z(P�M|)��L��*g7�2�2�WD��̐���8����Y���#����+��M.|��+�Ay���;����X�faE�o'^=�S��(�$�Z����B���>Ξ9��v����Ih����f�w�rS�3��[�2��` UUǢ>��GB\�m�zx����L�7l@f9��"M��_=�
hv�1Lr[��6  xt���7C��^݈�\b� E�Aj�4��ʨsy����.�S�z�8��oZ��Q����������#O����a}��~�o!����׺5$��Gb�K�����hk!���]�������� I���:��H�W�B��K^����>�eO����?�DKI��y�?I�m��x��� g�@'}I�	l����闁�H{�9�[^�<��V�5�c�C�T�����5/�Xi�3c�WU>�~��u�����[�����IE��I73��ZS�G�w/�+�i�y��u�p�"�E�N56�2��#�}�4 ��-�J��Ɵ~	{;��^>��X�?@��!_���|��@��B4�w�-�'�cm���B���+��HI��wD5:�.��
���7I�!Ϊ!N�Xԫ3�t��Xf�͖}�d��Xz��KHX��|Oˬ�� ��D	AHz������t?θ�ߣ�>h�\��A��<a'C(<A:ݏ����'	��	aj=���Q�N�~y�|`��'�-ޢ	��5�^���6�@���&U�ϕ]��JG�O<ѶwV��L�$8�����Q�ڂ������`g� '}	����̃krI}yH���i�Q�C�g\��27؏;ռ,�{oY �P/�������$���Q��1O�M*�*fi��7I_���Š�1(� g���-�!�;��ǻ7K���~��6�������|�c����m��B�� '
�~n��X��O����w��H��;�9 �'+�=>�y�+�'�d��0��`\�U�3���>v��#�õ�|��3f&��~��	�6��t����(����rT]Y����Q���O�ʁ1p�Z,�r8��t?ٸ��*A�D�G��/���S��!N��W��y����Z�����|̝���,i�x��W�a��h2��4=��߿?��ś���`0!����]�9;!�-���iC�J,M�MY�}����a�gk20C�������:���: �RvFH��:��eD�*�|��N�zV�dpP�I�,(�P�xKs�Sf%y�?I��-0=�"�!��4U�=u��w闥�ܣ��/���:;��	�Q�� ƫ!���U�V���e�Ɵ
��O󉦸��:��j�AS/(-���rJd�ui�c��>��Ԣ�IK�4;��	�;��j�zu�y���Nh���<�^��s�>] �������Yޞ6��V��D,{�$�"5
4@�~���p-�z(2�G�A�6�E^7re#
���)�ِ�6̹K1�O-�Hƫ94橇�����3{Z�@��޹@{⌵��]��.�2.��p>aҐ����aO��;��~�������̨6�~L��^2�*	�I��c DB#��Nb��^��(�j�\n�5Э�,�0n�S�qw����y5dǸ�/��GP'�W�&r��k��Լ�ϪE`/Aq�0 �_�'��c�Gu��:����'��%����r������8�u�br@���ׄ��@|/k��ƗRs�����)�;N!ۃ�x<��Q/_[�7��FB�@`�!W4������Mdm�Z���5���į��Җ��7�7Y(�99�(�= ҇���)3}�����y�vˑ��:��mN�觎����QT4��N;0�p�K�e�8-�m�Wf$�"�
�Z�K]E��/)Q������鰢I�_������P�W6��*%G�����Z0�������C��~����I��X��x3��tC���^�QCN�Eu^�_q���6�{��U"�2mxW-��og��p��750������ux	����O������Lwqeh�	��NT(����|���Y%��!��1&Ǫ����rp�t��m�=��/:&�\QXvg�AC�/��;����|��':�4�#�IT�i�J���w�0���f�N2>_��h1v�]�J¶�n�9M���{+	�[�#I/��c��X��a�4��$���c� [-�N�*������)B�Vf��Wn��aAg����֩O5. Eq��J.5��O����,'8�f��A)'ZX��U�	��
uƁX�F}�>�]��R�s��2w�7`�5�������/��>�ͣm4G7N	��$��x����w�`�e-��ܮ��<V2>��8]���f�vx���p��x��'ֶ�x�Ś�8���Q�9��w���i`>��iqH�/.���p8[�jVE1"�L����.�
U�(�O�B��u�����8��=�2][gb�����Xژ!?W�^jv~̰�;v�ŏ^�z9�''��-�sb2�[�;�VT��C�Ҙ���Bƚ��yq�MXU�u�����|(���ok�������y}b�Uv�׋�r�%�v�(_��eη�4�Ӷ��C��^4𕓬7\�D���r<r�,�p��Y<&��A�VS��V���]ay��wV�k۠��SI�?�l��3��	�5^��Z"����U^%��k4�/���q����q �}a}���%�ւ�߇�E�����ռ��c��v�S�M��|ׯ���9�`z�$2ѱs��|JJ�@0���K�H8�����|��#����x�OGó߮�G���4I���{��K�gX�?��~�1�_NmA��2�d�����c<�,-�x�7Qŀh/�}����u�A�y���)�K(���U0�V�#g�۪�ͧ�"�4�Gٯ`�����T��$+;��Z`S�Pw���		ko����Ys�<L��%X��ڗ� ����H�8ןA�
�/-���6�����oD@n�������7d�Lْ�ZJ��g�8� 6o%��ퟫ��fDq@2�KD�u�Q�]!0Fqz��x�Y �͓��f��I<|lw������_=��r���d��X�%�ق�r�Y�T�"<!�2���4�Q���������5�6�?�$�z�Ď\�ٮ, ����=������ ��T��u���5Ӥ���8`�fz���|�n���������7뀦��T�Ƥ��.�
��xsi���e���XB,�{R�t��5�o[���t�%h������I�cf��Fw���J��۲1P)�>�Y�X���Y�+� �.��m8��.��k$ߵ�����}�L�)�\��}{�����Qs�����J�(���I��׼��-��Пv�Ҫ��vPP8��Bv�`�Q��j^�!9P>B�6h�B )���%6gI��Ff8n����	�Ň�rii�����s���C�}�{��m\���K��+m��.�SB��L�ڵ�[��D����n��X6l���9��nO'����J�q1��\��F��CIy|~����)���4f��*衂�[��2��r�~u�|������;�ujy����Ǵ읕���/XDD����;U�+��_��n$�S���vv���T�����X"�O��鈬o�74�E_�V3����x66D�`���N�*��e�J���+1³7�dFe�O�K���Z��H��/�Ff��6��"�
j��\�*�bI �l>���o&����w��L�b��6�z>9�����00�#^�Kdґ��n_�:�ec�����ʲ��!�T���w��Q���]R��b����e?;�m�I(�������H��)�ikU�\�<)����t6x��l^T����0�u� 2B�G�_\�u�w	E�v�FD&�"�
Ƚ�H�V~�:�h<|�7���Bg�}S�L%fe��ܤ�L�p�_:�=#��J�x�&����ZL�ߌ'���B����W� E� 3*�ﭥz�M֛XQq� D
�7�r��0E�q����UJ����Z��<;OG!F��cVY��B&��f�n,N�B�ϣ��׳.��;����澸�7Y��v;�������O
M�L�^��)[e��1$����1�ra�G�i��*�])��Ns�2���e9:���C\�����ԅ=�+G2"w9r��F yUQ����p������?8�O�Hi؞�z*�_�b��&7���R~4�9O
(�_�� �L�!�6*�h�����h�g����?�ڶ J]�f����g�LO��v��{Si��@��OU����60DI�~H��\���I�u��^c�.�XM�L�$�qm��5w|�[m�6ak׸�R�}1����_Q{��������͌��2[y��-��J���&��f%[��b�N��7��R�N&I�.xH.E5� �����~�E�c�"*�ϩ����udcB�%B�U���Z�?�Z��5�Tj��4Ns8퉹��U�m(Qy�5,:��]��\lp���p�,gC0�amo�y��[ϰq�p��
/)g+􇙔��"�J֪%�gs�K��fKU�"���K�}�#�I������u�D]J��V�e���?�D�(�W9M�Q���Jq݄��vי	������\;��3>�Ə�
�w���U�G(��u���C����ׇ�V�r��(�e������0�3�B��AeU�|�g
E'��OL��_��F���=i\�ĝ$�[�hC�u�hM��KY�ڕui����J�Tie���V{�
�u)Bu%B�"�6~�U�:��r�|���}f��y�����m��Kk
�գ��B�~۾Գ!�fdk��4=��v"����9{�+��by�F}�l��x���C��.(��ܸ�
O�1ݚ������w�g�`�?+��Ƅ�����>�����bUb��!� ���QJ���[�q�Kb��[u��Vp#c�;z������+���W�����ͬ�S��_�±�"M�C��o������*0�sw� ���j�v�-����>yMg�n$��|⃸ti��S*i\��/���`��ڵ�=�����g�d1��]�˝��xU��&�MG��|�d�>�+}�ǃ���b�ya��̴5��%�˟�FR�n;E�#�v�3}��ݚJ��Lc5?��V�@�xP`����-<� �`WQ�x�S��xw�M��sA�FV��&�x;C �*�*�V׳9���p/\)��ƨ�)��#;���q�x��v��z�K�u�8�����I�u�׌����d$����z}�i��+{�ǁ��R{E~�F�5�@,�N4��i_�ǫ�о"�u|WR�dM�`�I���`$)�B�Ճ��t�\�^p�3y"+H�9τ��4�n�E���C������Upm�ѠQ��U����ifru$-���f�Y9o�g�,OKa��`����-��L[i�c���B�=�a����3�{6� ��p����+�r??,��=wh�z�c���L�Gf+u������A����zKP�C���A��Q��!��x��f�qX�5K�<���/o�0���85#�ԝ� �����S۞����8ɚ��u�-q��1h1Y����+$�c���V����^�d�E��Ñ�.�PI�!q�gԥ^����'�V'���#m*��NWC^��[��!��#F̙�;�w�$��mf@>�����y(���H�Q�U��*���Y�*�YԮ'L�t_q�yЯ^�,�Ɖ(��/�F���P��Q��3�m�䮹�o�}K

��*�uQ��2���+L��WN�A����0e���1�٬Z��"�cZ�n
J��g�R
�����F��B�����o�����\�XM��α�e�X;/��c��@���O8�ic��P���(�B��+;�ʗ�]7�T�u@*"oG��������s�\R^���̲-�8.��-L�GeT���R
�ˋ9Vs������Ŀ���:�d!�kJ�u��q�E0���.[�Y/��^/}��󮘾�R�ܓ��P�V�~u�?ö4��5A*���Ɍ�����<��Uhj�Y�;���*���)�c�X��1�U�����Z1g7�p��#�1��U:�C%�N��5�(�cȵ��񦰈?�ӭ�w�����������䵔.��p�h<��"(/u�(}��
G�g��T�[�I��H_��7�A��WlK���O��,*Vh_�Pih3}�7_�LM�t�hZĽo��)�-gI`��?O��W�Xf������^V���B����S��j�y,<5}�W ����'�Z��+�ψ@]KK��Ci�ۑZњM��/��*L�r�>���M S3�G����	����`d
��P�O�$��L� ���4�Ó�3�I@�.Α-S�2���i艶ͥ���F�T^Y�MtOL�+T#~�	�W�����!�P�;_�7��~���]��X���5p�"�>"��<�+����i �L_ظ�Bݬ2�v��ٳ�[�ޅ$�-��̬7���5X�~$�s�ʓ�C�����y���A�Fn�e��2����,JI6���.�
�t�Ø_�����0�5Zd��θ�����`����<�X�<�
PN�i�p_?�WK��~x��?�qO��7�P� �������oV��'��=�Ӯ��_����gDY��%�|��#��c� :sv�5���0�e7��F�%�|��kZ�)ʘ\�j}I;z��RvM� �eQi9�==�Ǌ�Zym�ˊ��g1gq�y@�3��c��t#�Ky� ��oٗ=0Mq�w�MY���ݩ��L9�"D�m�>3����[�~�8�,�M���^��Be=�	��'�~�8��F�D����}U��G�_�0>�(CJ�j�{�Ǯ��$��H�_)�V|����yo�,���ԩ�0fT��`J��w�	w�¹��u� ]:Q�뙏�ޛ�0�w��X�����|��k��	��%m�@��)�W��rnU�ӷ��¸��m��]���ev�8/��2��«ǰ����S�pK�
�q����f��>����%H!-G!�����/>��ok�M�xt�՝_�~K$j=(�PK   g�X�7}b  ]  /   images/89a9346c-9df8-41df-b8bd-ea49767937e0.png]��PNG

   IHDR   d   3   ai�   	pHYs  N�  N��"��   tEXtSoftware www.inkscape.org��<  �IDATx��\	��Wq����c�{gfgv��5۬/��)F���("�X�+R!"F�����#Aز�m6���]�w�;;;�s��3����w�����O���.�ݖ�7�]��zU��ޫ�^�]���>D��)wb�d�����p8J�M��x�Q��iH�xڇe�3̣��zI��V��ϝX&��\���U�9��:f��h�P���$X�pbf�!oV�+��
h������i&�j�fJ���Q��0��� �97:�bН%)���#F�w����<�%*�V'��z��fs��Qxg:f	��P
5�����i�Iöi���S�o0y�����)�C�����Q��7�{� 3���p��ӄQ�PG�!�U��;�a:�L��	̡�߻�s2�k�2�	�;�����8�eH�<J�Q�"ux�n�`DC&'��`�0\�`�5ޥ@z�, a_V�i�B�=����e����qd|l������E�{:ZW� ��E��{(Ң{��v!f�?Y�������)wsǌ#��q<?�B�%�*����М��B����ᖫV���qz�O�T���L	���&X��^ӖAS��'φ��u5���˵�^�:nqî$��������ݽ	��fI1�M}o��!�v�8�v ����XN�7���1�<�䲻����%0���ଯ���z�486v�3C3��SC!5��jΡ�)�Gτ�1)o���
�}��Q���Od�b�Nʏo`�)�ߦ�eXm�ؘ�.��ߝ$'��F�%�􌏤t=�����6�`��[	�$t"f@��D�If�ҷ���Й��I������^"WXc,!X%�6M#��(��"b�;+�$ac~�c[rK�J���.��?�u�|h38�X��k�R�f���1ˮ�W�c��^Ni&�X.�*نd�K�,AzYU�λK�D�E�
�'=�$uWI/�F�%�ؕ�`)��� ;Bm���:�t������7#}s���D���Ӥ�]�0���ۚ9ƶ��y��ʙbO�g1a��!�b��o�E��I.K+(�ؠ�P�pV"m�M�M�QOjP��2+o��l�4%@ӯ@_�`3�-�dn�k߇���Ͱj���c��H��drVJr4& �t���	�'�u;������Qlܽd���\T�E��P�D#�9�&"��^�	�6U=a��(ڝ��r�Rdx��!���(�</F4j�%�l�g���G��w��[xn��"�V�n�S���,X��1��V�4p���t�&Bv��P�,a��*	n3� �A�4�{�}���y�m�h�#�����(��wt�&Lj,����,����&��6"�/���4�B�p�:[���#3����Cس�C�?ta
��*Zښ���$��S���mGMM~�h`t|K�q�j/�~�&摜]$�;��gjk��,�p��d����#u����1��Z�;��X+}��� �UD��W��u#��`�ܸ_}C#:;��Leqfp��\�����	~�|���R�>�g%���㖲<�2C4|�8�
�Ģ�R%���l��M�%�]�o��d��	��H��Ko�V�5d`]N���ʩ���P���ġ���IֺX,PZ��2Lw�|����@*�&"9*�P���JR����&L����U�A��ԖN�x�j��`�}�v)U��_P�.]G.WRmҏ9T'���ߔ>G��K�_�Z��TFn�p�o�M��ot|Κ� �t*'F������
�h�Q��ф՚��XM��K�Ee�w��9�7=�$�`0�g���<�BmiV��Ό
���C��C�E ��@3��Bx�0>9O�Ε��Y���qJgrg!�2����2S�o�����ĩ��*��R�X���s?���VI�%$��a���vQ�]�Q�l��W~���tn�qc�[����L$�B���-x�bi���� �����N��l ;щELN/m��%1dc*)���'M-��1��b��084����;�N�q��I�����M��>���<�+�&Hsش��%uLل-�V+GL������XZZ�]w���_����'�p:���[m����xu���ɞ�������Z%�����u��O�63���"�m��������ӆ3���'n;�mm�HҶ�c��<r����|5�UV�|m�k�:9!�M/�gf�h�D[��ر��BKf���dd��%���<v6���r��Ѿ��ؠ�B~L�,���w|�3x��1ڳu��u�p���ٶ��,f
;����Rf��[*����,�y��7�=�N݃sS<��������*�F��jIL_�������S�s�\d���=�C��`�LY��>İ�&sCG�_�닸��G������|wC|��{��lY#������S��u̷��3��1C�]�Cf���&Ƹ���?��]�+9��7<C*��$�.�F2M�By��e��/��LF}��9����s�o?�.4ԇ�9��lr�Y?�啛��ێ��%�%Mՙ._U�,�6�ȯg��c�V|ʕSY�T�������(�JkOkR�07V��夻��V�; Q|�t۠�������(��ne�uy�:K~$�����o�:i	g1�⛿�AW�Mi<p��*a��.F�.�ZBg
z��x�/#\X������W/�POL���tgwCڒ���̹_uy�J3�
.�dc����ئU
۔]�)a'.[�����zJ�y��Sg�w�eqxw�4�//���L�d�t�^S�&u���C�꼁w����l�S�P�:����V���|܃唛�*�Huu��S_bWJ�oL��*��ģ���>�V�8�>O�������n��c��ӆ��9!�}��/h��c�rN��li�E׎f?y�޴�ӋXX\�C,���	��I������D"]�������*��thW� a5ľ�;n^�(#��K87�ώ��:� �O3����������o��_�^o�� �M ��������|��9O�L��_�w|���G߇��>bPZ��q�¤����j2#g���`����� O<����0�����<�����u�a2�����MfO�[ɠ��Z���S�g�3r�~����ŗ.���dp䅳��Ղw�z-j�|ph�iF}�� IG{[�̚���i�v2Y�ֆ09� G��\ՅPЏ=�;��{�M7�G��f^A�sYe�g�o�$����h�S7Y����5!>�|�]b+�6̱Cp�������VM��A�0��3���~�� >����} m��8sn���b��S������8���)L.�֫,���R*�Q��b�:1Ad)N�B�ňo؇G�|ѕU\����)Qao��]�z4�u�"���BLȡ���lC1켨���%��.3g��<Bjk�;���݊���T�V]���ZA�/���Gv�3��n��:ë�'|�$:k�djR�=�����f_�x��uV�RM��5�J;l+N�ˌ��3��y�lۈ���Ɍ`f2sy�����I�5��f����u�)�3���o�&vܵw6�=�p�/z�qg��n�^�sn;��XKj���;*�)֗S�e������Z��՗�Nx�{t�5����U�I�����:�d�{�� �E1�LM��e	6_�s_�.���W�L�h���λ������M*]'՜�����ǃ��O�^��
3!�+��<Fj�g�f�`��p�>��>���y��� ���7ϋ�2���5��͠���o	�xjU�d�����u��� �mwh��O�����+���]�;���j�q�����a"�W�Q�R��g���|a�[l�����L}n!Vv�t���k�z$���i�V$2.��mf��VY��Xd�*_T�\m^�jȞ@�&�~&�����m��28;p�--�����S����h)�yѠ���r�U��y+Icf��qo����=Q�U!�Wބ�ZKl�x���ބ��(b�8��owbp` �@ ���Sr�w���jo%��K5��J���ϊ��nI�
�3rE�kz�c]^��$/��Ey/��y11>�CC��|H�i	~��W���Č�]��юK��_cؐwv��ҒB�z%��.�PЇ��y���������;�W�]C����7�n��KM���'�����;W�0艧^Bm����rs��sϡ��7�r���En.^n��b�K�tPn���U�Ea���M��~�-�ު��iټ����M^�b	�������x\�`Ng+��pb�1�NDԫ�-�e<؁�#���'`��m�\N
��3rH�ʤv�k��H����񤱶��v��&5`Xul�z��Y�`��꟫���G�	&/������tխSG�o����m���6e����>�ۉ��4���G�mү�򂊗Y�)�B��+'Fpwo���W�i<w������߅��Z���3Y�85,������\�wp�.q�O�,b|rA}�v�s��%��oO'��=�L���:����?o��}t�h��؜<.�r�!�n/�i��>,���xF^4��r�Į��]��������s�s��ӄ���j���*F��RG��/Z	���=ޗF�u�^d�"��3gǅ��a|��ߧ�[��b�)�Q���(���y���~^eXXYB��Iĭ�|�`���I:�f��+�����D���-={�/,��cZ2�$lq9A,R{%�J*O3o��f��Nb�I��/�^���ȬH3�V�g
>�OpD���.��0F�%-m��T���r<��Ub�z�-�+���g��$p,�[̀{M�E�2�8'��-l3d�	����)�!7R�]�ɁD|	�ļ ����`bb���sI�K�4�#q!�a�h��[o��))ǁ���U���e5妁�H�F(�L@sx�r["6�Ċ������C,�����KF>���*�y���ޟk�o���22Ɉ�a�R��,]�*r!YD<�}����1��>L�1h,��g��D�dB�1ᮤ� �?GDP�+E��H����Vy���R���6n�yЛE{m\�ۨ�.ڿ$J	��9�連)��@$F] %Ag�eeM"�p���`w��8� �)�j���ql���0v�.��l܏�d������.�f��9ڄ��hJ`;ڄو��&8��S4T���`Rpb��,�֗�ߓ�%I``cZ+�E*M�m��J1ֳ�2�8��͕��fH�̢�;�Z�#����q�1b�	qdP�:�!W�Ys�S��80�S6��r�KĔ�Vua.+$�n�@H����J�S�7�'PD�`�DtuH��ƣ>�R�C��� �0��5��T.�х�!�R�M���c1�<u�nn=�Q(2���fB��pq8𘄧AL��Q|�.��7$<��R��M��� a��z�����k�۩�����o�|����l�WgZ�眛�єV����2¤�-�7KOc�.Y�rT9&�N��s�F�2��2��)<p�N��%?�1$��'�T�	�Wc&�N⡗k�-ZoΉ�o#�/�D@�0�����^��-3��p�R�f8�U�9�{_{�F��)���а�9+���p���b`+���ٰ�&�1��ud��S�"�<�0G,�MJt"���@~��^b����jl��J%C>C�����,TȠN�����D��χ�s(��[+�i�d�T���OPqY0V;cKLF��rr�鱁�2�$��	_y���-��,��c*���\PS����G��̡��0�ϯ΅����Ϗ��ݹ�h@چ�G<��S6��YqK@a�5�(1��ӢT��d���OBE`�G���Ǳ!�ɏ,6r���]f��$�ӎ���3D7s�2���G\k%�(G\sav���}������k�f�6����0�;Ov))1�x@���۰:�J���a�r�yC!϶��b�hk �dG���Nd֢ޑ�X*���^�.kE�c��ޱ�d|�g�D�c)ZQ�8��4{,�������L�����a#8�}�t�?��q�d�    IEND�B`�PK   k�X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   k�XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   ��X���  ~     jsons/user_defined.json���N�8�_���1���E�+�C3��i�F98�I�@����0��8S�W����q�/�O^�����U�5����(u,�G]7EU�h��؜i����_�l����m����=:��*I��i��۪~6�Ӳ�u�ۣ*?��+��&�Y!7oWm��EP��@�9�\�V�
�`:LRBC�B�XE�cBݤuqh�l?�-R�`E��y��!�(	U�P(��,Ͳ��塼5�iUڛ�	AY��*��M8��D&Y�c�Ddn��t��/�yXo���8����(O˼
V/A��o�氏����Y� �%��"3���E�4\3���Y�]�,:�T�iv��f�w����~V�����`��s>0�f]�wUmn~_�}��~���q8v������x��D�{��≃g�#(~w�S��{��	�_R/�9��Ν0�x�ܡKGL�^z���2\0��K]Yz��tJJ����3pN^���+�-��sr*屫Wl�	xy�Ο���,D��g����wE��F�g���?��[�.����ő]!毙��9�ગ0��R2�P��hxMS6U��/�|��|y�����c
���v5�{*��pE�B��̿m�v���S&��e���l.� ��+be� G��~����}xF�F� #�} A�	 �\c2,�f�� ��1^2��*q���U1�2�<��&�l�V��u<��#��daz�yJ���+kt�����Ws���n��Ҙ!iu�J]��w����ju�u�eut�=��qΊ����h�j�׵cp�&68B��3dl�(�a�Hʄ�3���'g$��g!M�
Y�U(y&B!t�SFx�7��?$=!�ϰ��UWV��)���1�b��<wb�����$���˓�-|��~ʅ�󋓿f��y@����#b��.�n��D�~�Hѓ 攊G
���P��k�N5nnA#���n	#|fN4h#���뉮��e�z�s%E`����_#��R�oYF\�RhA�
�c0b7�9 cv=U G:L`�I�5�)Pv�g���A�~!����C�~ю4�8�b��e����U�x	�N���Ɔ���j�	R'�+�a3�P'��ȾE��	C:�q1 u�l]H�����]��ټ��|���k@Q�;(	S�YȨ�Ä����INb�f��o�/�����Jc'jzh�!������Q������gk�����<6��ǌ{/�+�"���j����~y|����jcL~
m��=n��?��޼�PK
   ��X7���;!  )?                  cirkitFile.jsonPK
   g�X8�w���  ��  /             h!  images/219287a5-9258-450b-9fa3-793f4dcddf2e.pngPK
   g�X�7}b  ]  /             ��  images/89a9346c-9df8-41df-b8bd-ea49767937e0.pngPK
   k�X$7h�!  �!  /             c images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   k�XP��/�  ǽ  /             �/ images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   ��X���  ~               �� jsons/user_defined.jsonPK      �  9�   